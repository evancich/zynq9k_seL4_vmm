/*
 * Copyright 2017, Data61
 * Commonwealth Scientific and Industrial Research Organisation (CSIRO)
 * ABN 41 687 119 230.
 *
 * This software may be distributed and modified according to the terms of
 * the BSD 2-Clause license. Note that NO WARRANTY is provided.
 * See "LICENSE_BSD2.txt" for details.
 *
 * @TAG(DATA61_BSD)
 */

arch arm11

objects {
can_obj_7_0_control_9_tcb = tcb (addr: 0x13ae00, ip: 0x17848, sp: 0x14d000, elf: can_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [2], fault_ep: 0x00000003)
can_obj_7_0_fault_handler_15_0000_tcb = tcb (addr: 0x134e00, ip: 0x17848, sp: 0x141000, elf: can_obj_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [6])
can_obj_7_Int_3_0000_tcb = tcb (addr: 0x137e00, ip: 0x17848, sp: 0x147000, elf: can_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [4], fault_ep: 0x00000005)
can_obj_cnode = cnode (4 bits)
can_obj_fault_ep = ep
can_obj_group_bin_pd = pd
can_obj_interface_init_ep = ep
can_obj_m_test = notification
can_obj_post_init_ep = ep
can_obj_pre_init_ep = ep
can_spi_ep = ep
clk_obj_7_0_control_9_tcb = tcb (addr: 0x13ae00, ip: 0x14ce8, sp: 0x14d000, elf: clk_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [1], fault_ep: 0x00000002)
clk_obj_7_0_fault_handler_15_0000_tcb = tcb (addr: 0x134e00, ip: 0x14ce8, sp: 0x141000, elf: clk_obj_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [5])
clk_obj_7_clktree_7_0000_tcb = tcb (addr: 0x137e00, ip: 0x14ce8, sp: 0x147000, elf: clk_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [3], fault_ep: 0x00000004)
clk_obj_cnode = cnode (4 bits)
clk_obj_fault_ep = ep
clk_obj_group_bin_pd = pd
clk_obj_interface_init_ep = ep
clk_obj_post_init_ep = ep
clk_obj_pre_init_ep = ep
fd_pwm.vm_pwm_ep = ep
frame_can_obj_group_bin_0000 = frame (4k)
frame_can_obj_group_bin_0001 = frame (4k)
frame_can_obj_group_bin_0002 = frame (4k)
frame_can_obj_group_bin_0003 = frame (4k)
frame_can_obj_group_bin_0004 = frame (4k)
frame_can_obj_group_bin_0005 = frame (4k)
frame_can_obj_group_bin_0006 = frame (4k)
frame_can_obj_group_bin_0007 = frame (4k)
frame_can_obj_group_bin_0008 = frame (4k)
frame_can_obj_group_bin_0009 = frame (4k)
frame_can_obj_group_bin_0010 = frame (4k)
frame_can_obj_group_bin_0011 = frame (4k)
frame_can_obj_group_bin_0012 = frame (4k)
frame_can_obj_group_bin_0013 = frame (4k)
frame_can_obj_group_bin_0014 = frame (4k)
frame_can_obj_group_bin_0015 = frame (4k)
frame_can_obj_group_bin_0016 = frame (4k)
frame_can_obj_group_bin_0017 = frame (4k)
frame_can_obj_group_bin_0018 = frame (4k)
frame_can_obj_group_bin_0019 = frame (4k)
frame_can_obj_group_bin_0020 = frame (4k)
frame_can_obj_group_bin_0021 = frame (4k)
frame_can_obj_group_bin_0022 = frame (4k)
frame_can_obj_group_bin_0023 = frame (4k)
frame_can_obj_group_bin_0024 = frame (4k)
frame_can_obj_group_bin_0025 = frame (4k)
frame_can_obj_group_bin_0026 = frame (4k)
frame_can_obj_group_bin_0027 = frame (4k)
frame_can_obj_group_bin_0028 = frame (4k)
frame_can_obj_group_bin_0029 = frame (4k)
frame_can_obj_group_bin_0030 = frame (4k)
frame_can_obj_group_bin_0031 = frame (4k)
frame_can_obj_group_bin_0032 = frame (4k)
frame_can_obj_group_bin_0033 = frame (4k)
frame_can_obj_group_bin_0034 = frame (4k)
frame_can_obj_group_bin_0035 = frame (4k)
frame_can_obj_group_bin_0036 = frame (4k)
frame_can_obj_group_bin_0037 = frame (4k)
frame_can_obj_group_bin_0038 = frame (4k)
frame_can_obj_group_bin_0039 = frame (4k)
frame_can_obj_group_bin_0040 = frame (4k)
frame_can_obj_group_bin_0041 = frame (4k)
frame_can_obj_group_bin_0042 = frame (4k)
frame_can_obj_group_bin_0043 = frame (4k)
frame_can_obj_group_bin_0044 = frame (4k)
frame_can_obj_group_bin_0045 = frame (4k)
frame_can_obj_group_bin_0046 = frame (4k)
frame_can_obj_group_bin_0047 = frame (4k)
frame_can_obj_group_bin_0048 = frame (4k)
frame_can_obj_group_bin_0049 = frame (4k)
frame_can_obj_group_bin_0050 = frame (4k)
frame_can_obj_group_bin_0051 = frame (4k)
frame_can_obj_group_bin_0052 = frame (4k)
frame_can_obj_group_bin_0053 = frame (4k)
frame_can_obj_group_bin_0055 = frame (4k)
frame_can_obj_group_bin_0057 = frame (4k)
frame_can_obj_group_bin_0058 = frame (4k)
frame_can_obj_group_bin_0059 = frame (4k)
frame_can_obj_group_bin_0060 = frame (4k)
frame_can_obj_group_bin_0061 = frame (4k)
frame_can_obj_group_bin_0063 = frame (4k)
frame_can_obj_group_bin_0064 = frame (4k)
frame_can_obj_group_bin_0065 = frame (4k)
frame_can_obj_group_bin_0066 = frame (4k)
frame_can_obj_group_bin_0067 = frame (4k)
frame_can_obj_group_bin_0068 = frame (4k)
frame_can_obj_group_bin_0069 = frame (4k)
frame_can_obj_group_bin_0070 = frame (4k)
frame_can_obj_group_bin_0071 = frame (4k)
frame_can_obj_group_bin_0072 = frame (4k)
frame_can_obj_group_bin_0073 = frame (4k)
frame_can_obj_group_bin_0074 = frame (4k)
frame_can_obj_group_bin_0075 = frame (4k)
frame_can_obj_group_bin_0076 = frame (4k)
frame_can_obj_group_bin_0077 = frame (4k)
frame_can_obj_group_bin_0078 = frame (4k)
frame_can_obj_group_bin_0079 = frame (4k)
frame_can_obj_group_bin_0080 = frame (4k)
frame_can_obj_group_bin_0081 = frame (4k)
frame_can_obj_group_bin_0082 = frame (4k)
frame_can_obj_group_bin_0083 = frame (4k)
frame_can_obj_group_bin_0084 = frame (4k)
frame_can_obj_group_bin_0085 = frame (4k)
frame_can_obj_group_bin_0086 = frame (4k)
frame_can_obj_group_bin_0087 = frame (4k)
frame_can_obj_group_bin_0088 = frame (4k)
frame_can_obj_group_bin_0089 = frame (4k)
frame_can_obj_group_bin_0090 = frame (4k)
frame_can_obj_group_bin_0091 = frame (4k)
frame_can_obj_group_bin_0092 = frame (4k)
frame_can_obj_group_bin_0093 = frame (4k)
frame_can_obj_group_bin_0094 = frame (4k)
frame_can_obj_group_bin_0095 = frame (4k)
frame_can_obj_group_bin_0096 = frame (4k)
frame_can_obj_group_bin_0097 = frame (4k)
frame_can_obj_group_bin_0098 = frame (4k)
frame_can_obj_group_bin_0099 = frame (4k)
frame_can_obj_group_bin_0100 = frame (4k)
frame_can_obj_group_bin_0101 = frame (4k)
frame_can_obj_group_bin_0102 = frame (4k)
frame_can_obj_group_bin_0103 = frame (4k)
frame_can_obj_group_bin_0104 = frame (4k)
frame_can_obj_group_bin_0105 = frame (4k)
frame_can_obj_group_bin_0106 = frame (4k)
frame_can_obj_group_bin_0107 = frame (4k)
frame_can_obj_group_bin_0108 = frame (4k)
frame_can_obj_group_bin_0109 = frame (4k)
frame_can_obj_group_bin_0110 = frame (4k)
frame_can_obj_group_bin_0111 = frame (4k)
frame_can_obj_group_bin_0112 = frame (4k)
frame_can_obj_group_bin_0113 = frame (4k)
frame_can_obj_group_bin_0114 = frame (4k)
frame_can_obj_group_bin_0115 = frame (4k)
frame_can_obj_group_bin_0116 = frame (4k)
frame_can_obj_group_bin_0117 = frame (4k)
frame_can_obj_group_bin_0118 = frame (4k)
frame_can_obj_group_bin_0119 = frame (4k)
frame_can_obj_group_bin_0120 = frame (4k)
frame_can_obj_group_bin_0121 = frame (4k)
frame_can_obj_group_bin_0122 = frame (4k)
frame_can_obj_group_bin_0123 = frame (4k)
frame_can_obj_group_bin_0124 = frame (4k)
frame_can_obj_group_bin_0125 = frame (4k)
frame_can_obj_group_bin_0126 = frame (4k)
frame_can_obj_group_bin_0127 = frame (4k)
frame_can_obj_group_bin_0128 = frame (4k)
frame_can_obj_group_bin_0129 = frame (4k)
frame_can_obj_group_bin_0130 = frame (4k)
frame_can_obj_group_bin_0131 = frame (4k)
frame_can_obj_group_bin_0132 = frame (4k)
frame_can_obj_group_bin_0133 = frame (4k)
frame_can_obj_group_bin_0134 = frame (4k)
frame_can_obj_group_bin_0135 = frame (4k)
frame_can_obj_group_bin_0136 = frame (4k)
frame_can_obj_group_bin_0137 = frame (4k)
frame_can_obj_group_bin_0138 = frame (4k)
frame_can_obj_group_bin_0140 = frame (4k)
frame_can_obj_group_bin_0142 = frame (4k)
frame_can_obj_group_bin_0143 = frame (4k)
frame_can_obj_group_bin_0144 = frame (4k)
frame_can_obj_group_bin_0145 = frame (4k)
frame_can_obj_group_bin_0146 = frame (4k)
frame_can_obj_group_bin_0147 = frame (4k)
frame_can_obj_group_bin_0148 = frame (4k)
frame_can_obj_group_bin_0149 = frame (4k)
frame_can_obj_group_bin_0150 = frame (4k)
frame_can_obj_group_bin_0151 = frame (4k)
frame_can_obj_group_bin_0152 = frame (4k)
frame_can_obj_group_bin_0153 = frame (4k)
frame_can_obj_group_bin_0155 = frame (4k)
frame_can_obj_group_bin_0156 = frame (4k)
frame_can_obj_group_bin_0157 = frame (4k)
frame_can_obj_group_bin_0158 = frame (4k)
frame_can_obj_group_bin_0159 = frame (4k)
frame_can_obj_group_bin_0160 = frame (4k)
frame_can_obj_group_bin_0161 = frame (4k)
frame_can_obj_group_bin_0162 = frame (4k)
frame_can_obj_group_bin_0163 = frame (4k)
frame_can_obj_group_bin_0164 = frame (4k)
frame_can_obj_group_bin_0165 = frame (4k)
frame_can_obj_group_bin_0166 = frame (4k)
frame_can_obj_group_bin_0167 = frame (4k)
frame_can_obj_group_bin_0168 = frame (4k)
frame_can_obj_group_bin_0169 = frame (4k)
frame_can_obj_group_bin_0170 = frame (4k)
frame_can_obj_group_bin_0171 = frame (4k)
frame_can_obj_group_bin_0172 = frame (4k)
frame_can_obj_group_bin_0173 = frame (4k)
frame_can_obj_group_bin_0174 = frame (4k)
frame_can_obj_group_bin_0175 = frame (4k)
frame_can_obj_group_bin_0176 = frame (4k)
frame_can_obj_group_bin_0177 = frame (4k)
frame_can_obj_group_bin_0178 = frame (4k)
frame_can_obj_group_bin_0179 = frame (4k)
frame_can_obj_group_bin_0180 = frame (4k)
frame_can_obj_group_bin_0181 = frame (4k)
frame_can_obj_group_bin_0182 = frame (4k)
frame_can_obj_group_bin_0183 = frame (4k)
frame_can_obj_group_bin_0184 = frame (4k)
frame_can_obj_group_bin_0185 = frame (4k)
frame_can_obj_group_bin_0186 = frame (4k)
frame_can_obj_group_bin_0187 = frame (4k)
frame_can_obj_group_bin_0189 = frame (4k)
frame_can_obj_group_bin_0190 = frame (4k)
frame_can_obj_group_bin_0191 = frame (4k)
frame_can_obj_group_bin_0192 = frame (4k)
frame_can_obj_group_bin_0193 = frame (4k)
frame_can_obj_group_bin_0195 = frame (4k)
frame_can_obj_group_bin_0196 = frame (4k)
frame_can_obj_group_bin_0197 = frame (4k)
frame_can_obj_group_bin_0199 = frame (4k)
frame_can_obj_group_bin_0200 = frame (4k)
frame_can_obj_group_bin_0201 = frame (4k)
frame_can_obj_group_bin_0202 = frame (4k)
frame_can_obj_group_bin_0203 = frame (4k)
frame_can_obj_group_bin_0204 = frame (4k)
frame_can_obj_group_bin_0205 = frame (4k)
frame_can_obj_group_bin_0206 = frame (4k)
frame_can_obj_group_bin_0207 = frame (4k)
frame_can_obj_group_bin_0208 = frame (4k)
frame_can_obj_group_bin_0209 = frame (4k)
frame_can_obj_group_bin_0210 = frame (4k)
frame_can_obj_group_bin_0211 = frame (4k)
frame_can_obj_group_bin_0212 = frame (4k)
frame_can_obj_group_bin_0213 = frame (4k)
frame_can_obj_group_bin_0214 = frame (4k)
frame_can_obj_group_bin_0215 = frame (4k)
frame_can_obj_group_bin_0216 = frame (4k)
frame_can_obj_group_bin_0217 = frame (4k)
frame_can_obj_group_bin_0218 = frame (4k)
frame_can_obj_group_bin_0219 = frame (4k)
frame_can_obj_group_bin_0220 = frame (4k)
frame_can_obj_group_bin_0221 = frame (4k)
frame_can_obj_group_bin_0223 = frame (4k)
frame_can_obj_group_bin_0224 = frame (4k)
frame_can_obj_group_bin_0225 = frame (4k)
frame_can_obj_group_bin_0226 = frame (4k)
frame_can_obj_group_bin_0227 = frame (4k)
frame_can_obj_group_bin_0228 = frame (4k)
frame_can_obj_group_bin_0229 = frame (4k)
frame_can_obj_group_bin_0230 = frame (4k)
frame_can_obj_group_bin_0231 = frame (4k)
frame_can_obj_group_bin_0232 = frame (4k)
frame_can_obj_group_bin_0233 = frame (4k)
frame_can_obj_group_bin_0234 = frame (4k)
frame_can_obj_group_bin_0235 = frame (4k)
frame_can_obj_group_bin_0236 = frame (4k)
frame_can_obj_group_bin_0237 = frame (4k)
frame_can_obj_group_bin_0238 = frame (4k)
frame_can_obj_group_bin_0239 = frame (4k)
frame_can_obj_group_bin_0240 = frame (4k)
frame_can_obj_group_bin_0241 = frame (4k)
frame_can_obj_group_bin_0242 = frame (4k)
frame_can_obj_group_bin_0243 = frame (4k)
frame_can_obj_group_bin_0244 = frame (4k)
frame_can_obj_group_bin_0245 = frame (4k)
frame_can_obj_group_bin_0246 = frame (4k)
frame_can_obj_group_bin_0247 = frame (4k)
frame_can_obj_group_bin_0248 = frame (4k)
frame_can_obj_group_bin_0249 = frame (4k)
frame_can_obj_group_bin_0250 = frame (4k)
frame_can_obj_group_bin_0251 = frame (4k)
frame_can_obj_group_bin_0252 = frame (4k)
frame_can_obj_group_bin_0253 = frame (4k)
frame_can_obj_group_bin_0254 = frame (4k)
frame_can_obj_group_bin_0255 = frame (4k)
frame_can_obj_group_bin_0256 = frame (4k)
frame_can_obj_group_bin_0257 = frame (4k)
frame_can_obj_group_bin_0258 = frame (4k)
frame_can_obj_group_bin_0260 = frame (4k)
frame_can_obj_group_bin_0261 = frame (4k)
frame_can_obj_group_bin_0262 = frame (4k)
frame_can_obj_group_bin_0263 = frame (4k)
frame_can_obj_group_bin_0264 = frame (4k)
frame_can_obj_group_bin_0265 = frame (4k)
frame_can_obj_group_bin_0266 = frame (4k)
frame_can_obj_group_bin_0267 = frame (4k)
frame_can_obj_group_bin_0268 = frame (4k)
frame_can_obj_group_bin_0269 = frame (4k)
frame_can_obj_group_bin_0270 = frame (4k)
frame_can_obj_group_bin_0271 = frame (4k)
frame_can_obj_group_bin_0272 = frame (4k)
frame_can_obj_group_bin_0273 = frame (4k)
frame_can_obj_group_bin_0274 = frame (4k)
frame_can_obj_group_bin_0275 = frame (4k)
frame_can_obj_group_bin_0276 = frame (4k)
frame_can_obj_group_bin_0277 = frame (4k)
frame_can_obj_group_bin_0279 = frame (4k)
frame_can_obj_group_bin_0280 = frame (4k)
frame_can_obj_group_bin_0281 = frame (4k)
frame_can_obj_group_bin_0282 = frame (4k)
frame_can_obj_group_bin_0283 = frame (4k)
frame_can_obj_group_bin_0284 = frame (4k)
frame_can_obj_group_bin_0285 = frame (4k)
frame_can_obj_group_bin_0286 = frame (4k)
frame_can_obj_group_bin_0287 = frame (4k)
frame_can_obj_group_bin_0288 = frame (4k)
frame_can_obj_group_bin_0289 = frame (4k)
frame_can_obj_group_bin_0290 = frame (4k)
frame_can_obj_group_bin_0291 = frame (4k)
frame_can_obj_group_bin_0292 = frame (4k)
frame_can_obj_group_bin_0293 = frame (4k)
frame_can_obj_group_bin_0294 = frame (4k)
frame_can_obj_group_bin_0295 = frame (4k)
frame_can_obj_group_bin_0296 = frame (4k)
frame_can_obj_group_bin_0297 = frame (4k)
frame_can_obj_group_bin_0298 = frame (4k)
frame_can_obj_group_bin_0299 = frame (4k)
frame_can_obj_group_bin_0300 = frame (4k)
frame_can_obj_group_bin_0301 = frame (4k)
frame_can_obj_group_bin_0302 = frame (4k)
frame_can_obj_group_bin_0303 = frame (4k)
frame_clk_obj_group_bin_0000 = frame (4k)
frame_clk_obj_group_bin_0001 = frame (4k)
frame_clk_obj_group_bin_0002 = frame (4k)
frame_clk_obj_group_bin_0003 = frame (4k)
frame_clk_obj_group_bin_0004 = frame (4k)
frame_clk_obj_group_bin_0005 = frame (4k)
frame_clk_obj_group_bin_0006 = frame (4k)
frame_clk_obj_group_bin_0007 = frame (4k)
frame_clk_obj_group_bin_0008 = frame (4k)
frame_clk_obj_group_bin_0009 = frame (4k)
frame_clk_obj_group_bin_0010 = frame (4k)
frame_clk_obj_group_bin_0011 = frame (4k)
frame_clk_obj_group_bin_0012 = frame (4k)
frame_clk_obj_group_bin_0013 = frame (4k)
frame_clk_obj_group_bin_0014 = frame (4k)
frame_clk_obj_group_bin_0015 = frame (4k)
frame_clk_obj_group_bin_0016 = frame (4k)
frame_clk_obj_group_bin_0017 = frame (4k)
frame_clk_obj_group_bin_0018 = frame (4k)
frame_clk_obj_group_bin_0019 = frame (4k)
frame_clk_obj_group_bin_0020 = frame (4k)
frame_clk_obj_group_bin_0021 = frame (4k)
frame_clk_obj_group_bin_0022 = frame (4k)
frame_clk_obj_group_bin_0023 = frame (4k)
frame_clk_obj_group_bin_0024 = frame (4k)
frame_clk_obj_group_bin_0025 = frame (4k)
frame_clk_obj_group_bin_0026 = frame (4k)
frame_clk_obj_group_bin_0027 = frame (4k)
frame_clk_obj_group_bin_0028 = frame (4k)
frame_clk_obj_group_bin_0029 = frame (4k)
frame_clk_obj_group_bin_0030 = frame (4k)
frame_clk_obj_group_bin_0031 = frame (4k)
frame_clk_obj_group_bin_0032 = frame (4k)
frame_clk_obj_group_bin_0033 = frame (4k)
frame_clk_obj_group_bin_0034 = frame (4k)
frame_clk_obj_group_bin_0035 = frame (4k)
frame_clk_obj_group_bin_0036 = frame (4k)
frame_clk_obj_group_bin_0037 = frame (4k)
frame_clk_obj_group_bin_0038 = frame (4k)
frame_clk_obj_group_bin_0039 = frame (4k)
frame_clk_obj_group_bin_0040 = frame (4k)
frame_clk_obj_group_bin_0041 = frame (4k)
frame_clk_obj_group_bin_0042 = frame (4k)
frame_clk_obj_group_bin_0043 = frame (4k)
frame_clk_obj_group_bin_0044 = frame (4k)
frame_clk_obj_group_bin_0045 = frame (4k)
frame_clk_obj_group_bin_0046 = frame (4k)
frame_clk_obj_group_bin_0047 = frame (4k)
frame_clk_obj_group_bin_0048 = frame (4k)
frame_clk_obj_group_bin_0049 = frame (4k)
frame_clk_obj_group_bin_0050 = frame (4k)
frame_clk_obj_group_bin_0051 = frame (4k)
frame_clk_obj_group_bin_0052 = frame (4k)
frame_clk_obj_group_bin_0053 = frame (4k)
frame_clk_obj_group_bin_0055 = frame (4k)
frame_clk_obj_group_bin_0057 = frame (4k)
frame_clk_obj_group_bin_0058 = frame (4k)
frame_clk_obj_group_bin_0059 = frame (4k)
frame_clk_obj_group_bin_0060 = frame (4k)
frame_clk_obj_group_bin_0061 = frame (4k)
frame_clk_obj_group_bin_0063 = frame (4k)
frame_clk_obj_group_bin_0064 = frame (4k)
frame_clk_obj_group_bin_0065 = frame (4k)
frame_clk_obj_group_bin_0066 = frame (4k)
frame_clk_obj_group_bin_0067 = frame (4k)
frame_clk_obj_group_bin_0068 = frame (4k)
frame_clk_obj_group_bin_0069 = frame (4k)
frame_clk_obj_group_bin_0070 = frame (4k)
frame_clk_obj_group_bin_0071 = frame (4k)
frame_clk_obj_group_bin_0072 = frame (4k)
frame_clk_obj_group_bin_0073 = frame (4k)
frame_clk_obj_group_bin_0074 = frame (4k)
frame_clk_obj_group_bin_0075 = frame (4k)
frame_clk_obj_group_bin_0076 = frame (4k)
frame_clk_obj_group_bin_0077 = frame (4k)
frame_clk_obj_group_bin_0078 = frame (4k)
frame_clk_obj_group_bin_0079 = frame (4k)
frame_clk_obj_group_bin_0080 = frame (4k)
frame_clk_obj_group_bin_0081 = frame (4k)
frame_clk_obj_group_bin_0082 = frame (4k)
frame_clk_obj_group_bin_0083 = frame (4k)
frame_clk_obj_group_bin_0084 = frame (4k)
frame_clk_obj_group_bin_0085 = frame (4k)
frame_clk_obj_group_bin_0086 = frame (4k)
frame_clk_obj_group_bin_0087 = frame (4k)
frame_clk_obj_group_bin_0088 = frame (4k)
frame_clk_obj_group_bin_0089 = frame (4k)
frame_clk_obj_group_bin_0090 = frame (4k)
frame_clk_obj_group_bin_0091 = frame (4k)
frame_clk_obj_group_bin_0092 = frame (4k)
frame_clk_obj_group_bin_0093 = frame (4k)
frame_clk_obj_group_bin_0094 = frame (4k)
frame_clk_obj_group_bin_0095 = frame (4k)
frame_clk_obj_group_bin_0096 = frame (4k)
frame_clk_obj_group_bin_0097 = frame (4k)
frame_clk_obj_group_bin_0098 = frame (4k)
frame_clk_obj_group_bin_0099 = frame (4k)
frame_clk_obj_group_bin_0100 = frame (4k)
frame_clk_obj_group_bin_0101 = frame (4k)
frame_clk_obj_group_bin_0102 = frame (4k)
frame_clk_obj_group_bin_0103 = frame (4k)
frame_clk_obj_group_bin_0104 = frame (4k)
frame_clk_obj_group_bin_0105 = frame (4k, paddr: 0x10020000)
frame_clk_obj_group_bin_0106 = frame (4k)
frame_clk_obj_group_bin_0107 = frame (4k)
frame_clk_obj_group_bin_0108 = frame (4k)
frame_clk_obj_group_bin_0109 = frame (4k)
frame_clk_obj_group_bin_0110 = frame (4k)
frame_clk_obj_group_bin_0111 = frame (4k)
frame_clk_obj_group_bin_0112 = frame (4k)
frame_clk_obj_group_bin_0113 = frame (4k)
frame_clk_obj_group_bin_0114 = frame (4k)
frame_clk_obj_group_bin_0115 = frame (4k)
frame_clk_obj_group_bin_0116 = frame (4k)
frame_clk_obj_group_bin_0117 = frame (4k)
frame_clk_obj_group_bin_0118 = frame (4k)
frame_clk_obj_group_bin_0119 = frame (4k)
frame_clk_obj_group_bin_0120 = frame (4k)
frame_clk_obj_group_bin_0121 = frame (4k)
frame_clk_obj_group_bin_0122 = frame (4k)
frame_clk_obj_group_bin_0123 = frame (4k)
frame_clk_obj_group_bin_0124 = frame (4k)
frame_clk_obj_group_bin_0125 = frame (4k)
frame_clk_obj_group_bin_0126 = frame (4k)
frame_clk_obj_group_bin_0127 = frame (4k)
frame_clk_obj_group_bin_0128 = frame (4k)
frame_clk_obj_group_bin_0129 = frame (4k)
frame_clk_obj_group_bin_0130 = frame (4k)
frame_clk_obj_group_bin_0131 = frame (4k)
frame_clk_obj_group_bin_0132 = frame (4k)
frame_clk_obj_group_bin_0133 = frame (4k)
frame_clk_obj_group_bin_0134 = frame (4k)
frame_clk_obj_group_bin_0135 = frame (4k)
frame_clk_obj_group_bin_0136 = frame (4k)
frame_clk_obj_group_bin_0137 = frame (4k)
frame_clk_obj_group_bin_0138 = frame (4k)
frame_clk_obj_group_bin_0139 = frame (4k)
frame_clk_obj_group_bin_0141 = frame (4k)
frame_clk_obj_group_bin_0143 = frame (4k)
frame_clk_obj_group_bin_0144 = frame (4k)
frame_clk_obj_group_bin_0145 = frame (4k)
frame_clk_obj_group_bin_0146 = frame (4k)
frame_clk_obj_group_bin_0147 = frame (4k)
frame_clk_obj_group_bin_0148 = frame (4k)
frame_clk_obj_group_bin_0149 = frame (4k)
frame_clk_obj_group_bin_0150 = frame (4k)
frame_clk_obj_group_bin_0151 = frame (4k)
frame_clk_obj_group_bin_0152 = frame (4k)
frame_clk_obj_group_bin_0153 = frame (4k)
frame_clk_obj_group_bin_0154 = frame (4k)
frame_clk_obj_group_bin_0156 = frame (4k)
frame_clk_obj_group_bin_0157 = frame (4k)
frame_clk_obj_group_bin_0158 = frame (4k)
frame_clk_obj_group_bin_0159 = frame (4k)
frame_clk_obj_group_bin_0160 = frame (4k)
frame_clk_obj_group_bin_0161 = frame (4k)
frame_clk_obj_group_bin_0162 = frame (4k)
frame_clk_obj_group_bin_0163 = frame (4k)
frame_clk_obj_group_bin_0164 = frame (4k)
frame_clk_obj_group_bin_0165 = frame (4k)
frame_clk_obj_group_bin_0166 = frame (4k)
frame_clk_obj_group_bin_0167 = frame (4k)
frame_clk_obj_group_bin_0168 = frame (4k)
frame_clk_obj_group_bin_0169 = frame (4k)
frame_clk_obj_group_bin_0170 = frame (4k)
frame_clk_obj_group_bin_0171 = frame (4k)
frame_clk_obj_group_bin_0172 = frame (4k)
frame_clk_obj_group_bin_0173 = frame (4k)
frame_clk_obj_group_bin_0174 = frame (4k)
frame_clk_obj_group_bin_0175 = frame (4k)
frame_clk_obj_group_bin_0176 = frame (4k)
frame_clk_obj_group_bin_0177 = frame (4k)
frame_clk_obj_group_bin_0178 = frame (4k)
frame_clk_obj_group_bin_0179 = frame (4k)
frame_clk_obj_group_bin_0180 = frame (4k)
frame_clk_obj_group_bin_0181 = frame (4k)
frame_clk_obj_group_bin_0182 = frame (4k)
frame_clk_obj_group_bin_0183 = frame (4k)
frame_clk_obj_group_bin_0184 = frame (4k)
frame_clk_obj_group_bin_0185 = frame (4k)
frame_clk_obj_group_bin_0186 = frame (4k)
frame_clk_obj_group_bin_0187 = frame (4k)
frame_clk_obj_group_bin_0188 = frame (4k)
frame_clk_obj_group_bin_0190 = frame (4k)
frame_clk_obj_group_bin_0191 = frame (4k)
frame_clk_obj_group_bin_0192 = frame (4k)
frame_clk_obj_group_bin_0193 = frame (4k)
frame_clk_obj_group_bin_0194 = frame (4k)
frame_clk_obj_group_bin_0196 = frame (4k)
frame_clk_obj_group_bin_0197 = frame (4k)
frame_clk_obj_group_bin_0198 = frame (4k)
frame_clk_obj_group_bin_0200 = frame (4k)
frame_clk_obj_group_bin_0201 = frame (4k)
frame_clk_obj_group_bin_0202 = frame (4k)
frame_clk_obj_group_bin_0203 = frame (4k)
frame_clk_obj_group_bin_0204 = frame (4k)
frame_clk_obj_group_bin_0205 = frame (4k)
frame_clk_obj_group_bin_0206 = frame (4k)
frame_clk_obj_group_bin_0207 = frame (4k)
frame_clk_obj_group_bin_0208 = frame (4k)
frame_clk_obj_group_bin_0209 = frame (4k)
frame_clk_obj_group_bin_0210 = frame (4k)
frame_clk_obj_group_bin_0211 = frame (4k)
frame_clk_obj_group_bin_0212 = frame (4k)
frame_clk_obj_group_bin_0213 = frame (4k)
frame_clk_obj_group_bin_0214 = frame (4k)
frame_clk_obj_group_bin_0215 = frame (4k)
frame_clk_obj_group_bin_0216 = frame (4k)
frame_clk_obj_group_bin_0217 = frame (4k)
frame_clk_obj_group_bin_0218 = frame (4k)
frame_clk_obj_group_bin_0219 = frame (4k)
frame_clk_obj_group_bin_0220 = frame (4k)
frame_clk_obj_group_bin_0221 = frame (4k)
frame_clk_obj_group_bin_0222 = frame (4k)
frame_clk_obj_group_bin_0224 = frame (4k)
frame_clk_obj_group_bin_0225 = frame (4k)
frame_clk_obj_group_bin_0226 = frame (4k)
frame_clk_obj_group_bin_0227 = frame (4k)
frame_clk_obj_group_bin_0228 = frame (4k)
frame_clk_obj_group_bin_0229 = frame (4k)
frame_clk_obj_group_bin_0230 = frame (4k)
frame_clk_obj_group_bin_0231 = frame (4k)
frame_clk_obj_group_bin_0232 = frame (4k)
frame_clk_obj_group_bin_0233 = frame (4k)
frame_clk_obj_group_bin_0234 = frame (4k)
frame_clk_obj_group_bin_0235 = frame (4k)
frame_clk_obj_group_bin_0236 = frame (4k)
frame_clk_obj_group_bin_0237 = frame (4k)
frame_clk_obj_group_bin_0238 = frame (4k)
frame_clk_obj_group_bin_0239 = frame (4k, paddr: 0x10010000)
frame_clk_obj_group_bin_0240 = frame (4k)
frame_clk_obj_group_bin_0241 = frame (4k)
frame_clk_obj_group_bin_0242 = frame (4k)
frame_clk_obj_group_bin_0243 = frame (4k)
frame_clk_obj_group_bin_0244 = frame (4k)
frame_clk_obj_group_bin_0245 = frame (4k)
frame_clk_obj_group_bin_0246 = frame (4k)
frame_clk_obj_group_bin_0247 = frame (4k)
frame_clk_obj_group_bin_0248 = frame (4k)
frame_clk_obj_group_bin_0249 = frame (4k)
frame_clk_obj_group_bin_0250 = frame (4k)
frame_clk_obj_group_bin_0251 = frame (4k)
frame_clk_obj_group_bin_0252 = frame (4k)
frame_clk_obj_group_bin_0253 = frame (4k)
frame_clk_obj_group_bin_0254 = frame (4k)
frame_clk_obj_group_bin_0255 = frame (4k)
frame_clk_obj_group_bin_0256 = frame (4k)
frame_clk_obj_group_bin_0257 = frame (4k)
frame_clk_obj_group_bin_0258 = frame (4k)
frame_clk_obj_group_bin_0259 = frame (4k)
frame_clk_obj_group_bin_0260 = frame (4k)
frame_clk_obj_group_bin_0262 = frame (4k)
frame_clk_obj_group_bin_0263 = frame (4k)
frame_clk_obj_group_bin_0264 = frame (4k)
frame_clk_obj_group_bin_0265 = frame (4k)
frame_clk_obj_group_bin_0266 = frame (4k)
frame_clk_obj_group_bin_0267 = frame (4k)
frame_clk_obj_group_bin_0268 = frame (4k)
frame_clk_obj_group_bin_0269 = frame (4k)
frame_clk_obj_group_bin_0270 = frame (4k)
frame_clk_obj_group_bin_0271 = frame (4k)
frame_clk_obj_group_bin_0272 = frame (4k)
frame_clk_obj_group_bin_0273 = frame (4k)
frame_clk_obj_group_bin_0274 = frame (4k)
frame_clk_obj_group_bin_0275 = frame (4k)
frame_clk_obj_group_bin_0276 = frame (4k)
frame_clk_obj_group_bin_0277 = frame (4k)
frame_clk_obj_group_bin_0278 = frame (4k)
frame_clk_obj_group_bin_0279 = frame (4k)
frame_clk_obj_group_bin_0281 = frame (4k)
frame_clk_obj_group_bin_0282 = frame (4k)
frame_clk_obj_group_bin_0283 = frame (4k, paddr: 0x10014000)
frame_clk_obj_group_bin_0284 = frame (4k)
frame_clk_obj_group_bin_0285 = frame (4k)
frame_clk_obj_group_bin_0286 = frame (4k)
frame_clk_obj_group_bin_0287 = frame (4k)
frame_clk_obj_group_bin_0288 = frame (4k)
frame_clk_obj_group_bin_0289 = frame (4k)
frame_clk_obj_group_bin_0290 = frame (4k)
frame_clk_obj_group_bin_0291 = frame (4k)
frame_clk_obj_group_bin_0292 = frame (4k)
frame_clk_obj_group_bin_0293 = frame (4k)
frame_clk_obj_group_bin_0294 = frame (4k)
frame_clk_obj_group_bin_0295 = frame (4k)
frame_clk_obj_group_bin_0296 = frame (4k)
frame_clk_obj_group_bin_0297 = frame (4k)
frame_clk_obj_group_bin_0298 = frame (4k)
frame_clk_obj_group_bin_0299 = frame (4k)
frame_clk_obj_group_bin_0300 = frame (4k)
frame_clk_obj_group_bin_0301 = frame (4k)
frame_clk_obj_group_bin_0302 = frame (4k)
frame_clk_obj_group_bin_0303 = frame (4k)
frame_clk_obj_group_bin_0304 = frame (4k)
frame_clk_obj_group_bin_0305 = frame (4k)
frame_gpio_obj_group_bin_0000 = frame (4k)
frame_gpio_obj_group_bin_0001 = frame (4k)
frame_gpio_obj_group_bin_0002 = frame (4k)
frame_gpio_obj_group_bin_0003 = frame (4k)
frame_gpio_obj_group_bin_0004 = frame (4k)
frame_gpio_obj_group_bin_0005 = frame (4k)
frame_gpio_obj_group_bin_0006 = frame (4k, paddr: 0x13400000)
frame_gpio_obj_group_bin_0008 = frame (4k)
frame_gpio_obj_group_bin_0009 = frame (4k)
frame_gpio_obj_group_bin_0010 = frame (4k)
frame_gpio_obj_group_bin_0011 = frame (4k)
frame_gpio_obj_group_bin_0012 = frame (4k)
frame_gpio_obj_group_bin_0013 = frame (4k)
frame_gpio_obj_group_bin_0014 = frame (4k)
frame_gpio_obj_group_bin_0015 = frame (4k)
frame_gpio_obj_group_bin_0017 = frame (4k)
frame_gpio_obj_group_bin_0018 = frame (4k)
frame_gpio_obj_group_bin_0019 = frame (4k)
frame_gpio_obj_group_bin_0020 = frame (4k)
frame_gpio_obj_group_bin_0021 = frame (4k)
frame_gpio_obj_group_bin_0022 = frame (4k)
frame_gpio_obj_group_bin_0023 = frame (4k)
frame_gpio_obj_group_bin_0024 = frame (4k)
frame_gpio_obj_group_bin_0025 = frame (4k)
frame_gpio_obj_group_bin_0026 = frame (4k)
frame_gpio_obj_group_bin_0027 = frame (4k)
frame_gpio_obj_group_bin_0028 = frame (4k)
frame_gpio_obj_group_bin_0029 = frame (4k)
frame_gpio_obj_group_bin_0030 = frame (4k)
frame_gpio_obj_group_bin_0031 = frame (4k)
frame_gpio_obj_group_bin_0032 = frame (4k)
frame_gpio_obj_group_bin_0033 = frame (4k)
frame_gpio_obj_group_bin_0035 = frame (4k)
frame_gpio_obj_group_bin_0036 = frame (4k)
frame_gpio_obj_group_bin_0037 = frame (4k)
frame_gpio_obj_group_bin_0038 = frame (4k)
frame_gpio_obj_group_bin_0039 = frame (4k)
frame_gpio_obj_group_bin_0040 = frame (4k)
frame_gpio_obj_group_bin_0041 = frame (4k)
frame_gpio_obj_group_bin_0042 = frame (4k)
frame_gpio_obj_group_bin_0043 = frame (4k)
frame_gpio_obj_group_bin_0044 = frame (4k)
frame_gpio_obj_group_bin_0046 = frame (4k)
frame_gpio_obj_group_bin_0047 = frame (4k)
frame_gpio_obj_group_bin_0049 = frame (4k)
frame_gpio_obj_group_bin_0050 = frame (4k, paddr: 0x10440000)
frame_gpio_obj_group_bin_0051 = frame (4k)
frame_gpio_obj_group_bin_0052 = frame (4k)
frame_gpio_obj_group_bin_0053 = frame (4k)
frame_gpio_obj_group_bin_0054 = frame (4k)
frame_gpio_obj_group_bin_0055 = frame (4k)
frame_gpio_obj_group_bin_0057 = frame (4k)
frame_gpio_obj_group_bin_0058 = frame (4k)
frame_gpio_obj_group_bin_0059 = frame (4k)
frame_gpio_obj_group_bin_0060 = frame (4k)
frame_gpio_obj_group_bin_0061 = frame (4k)
frame_gpio_obj_group_bin_0062 = frame (4k)
frame_gpio_obj_group_bin_0063 = frame (4k)
frame_gpio_obj_group_bin_0064 = frame (4k)
frame_gpio_obj_group_bin_0065 = frame (4k)
frame_gpio_obj_group_bin_0066 = frame (4k)
frame_gpio_obj_group_bin_0067 = frame (4k)
frame_gpio_obj_group_bin_0068 = frame (4k)
frame_gpio_obj_group_bin_0069 = frame (4k)
frame_gpio_obj_group_bin_0070 = frame (4k)
frame_gpio_obj_group_bin_0071 = frame (4k)
frame_gpio_obj_group_bin_0072 = frame (4k)
frame_gpio_obj_group_bin_0073 = frame (4k)
frame_gpio_obj_group_bin_0074 = frame (4k)
frame_gpio_obj_group_bin_0075 = frame (4k)
frame_gpio_obj_group_bin_0076 = frame (4k)
frame_gpio_obj_group_bin_0078 = frame (4k)
frame_gpio_obj_group_bin_0079 = frame (4k)
frame_gpio_obj_group_bin_0080 = frame (4k)
frame_gpio_obj_group_bin_0081 = frame (4k)
frame_gpio_obj_group_bin_0082 = frame (4k)
frame_gpio_obj_group_bin_0083 = frame (4k)
frame_gpio_obj_group_bin_0084 = frame (4k)
frame_gpio_obj_group_bin_0085 = frame (4k)
frame_gpio_obj_group_bin_0086 = frame (4k)
frame_gpio_obj_group_bin_0088 = frame (4k)
frame_gpio_obj_group_bin_0089 = frame (4k)
frame_gpio_obj_group_bin_0091 = frame (4k)
frame_gpio_obj_group_bin_0092 = frame (4k)
frame_gpio_obj_group_bin_0093 = frame (4k)
frame_gpio_obj_group_bin_0094 = frame (4k)
frame_gpio_obj_group_bin_0096 = frame (4k)
frame_gpio_obj_group_bin_0097 = frame (4k)
frame_gpio_obj_group_bin_0098 = frame (4k)
frame_gpio_obj_group_bin_0099 = frame (4k)
frame_gpio_obj_group_bin_0100 = frame (4k)
frame_gpio_obj_group_bin_0101 = frame (4k)
frame_gpio_obj_group_bin_0102 = frame (4k)
frame_gpio_obj_group_bin_0103 = frame (4k)
frame_gpio_obj_group_bin_0104 = frame (4k)
frame_gpio_obj_group_bin_0105 = frame (4k)
frame_gpio_obj_group_bin_0106 = frame (4k)
frame_gpio_obj_group_bin_0107 = frame (4k)
frame_gpio_obj_group_bin_0108 = frame (4k)
frame_gpio_obj_group_bin_0109 = frame (4k)
frame_gpio_obj_group_bin_0110 = frame (4k)
frame_gpio_obj_group_bin_0111 = frame (4k)
frame_gpio_obj_group_bin_0112 = frame (4k)
frame_gpio_obj_group_bin_0113 = frame (4k)
frame_gpio_obj_group_bin_0114 = frame (4k)
frame_gpio_obj_group_bin_0115 = frame (4k)
frame_gpio_obj_group_bin_0117 = frame (4k)
frame_gpio_obj_group_bin_0118 = frame (4k)
frame_gpio_obj_group_bin_0119 = frame (4k)
frame_gpio_obj_group_bin_0120 = frame (4k)
frame_gpio_obj_group_bin_0121 = frame (4k)
frame_gpio_obj_group_bin_0122 = frame (4k)
frame_gpio_obj_group_bin_0123 = frame (4k)
frame_gpio_obj_group_bin_0124 = frame (4k)
frame_gpio_obj_group_bin_0125 = frame (4k)
frame_gpio_obj_group_bin_0126 = frame (4k)
frame_gpio_obj_group_bin_0128 = frame (4k)
frame_gpio_obj_group_bin_0130 = frame (4k)
frame_gpio_obj_group_bin_0131 = frame (4k)
frame_gpio_obj_group_bin_0132 = frame (4k)
frame_gpio_obj_group_bin_0133 = frame (4k)
frame_gpio_obj_group_bin_0134 = frame (4k)
frame_gpio_obj_group_bin_0135 = frame (4k)
frame_gpio_obj_group_bin_0136 = frame (4k)
frame_gpio_obj_group_bin_0138 = frame (4k)
frame_gpio_obj_group_bin_0139 = frame (4k)
frame_gpio_obj_group_bin_0140 = frame (4k)
frame_gpio_obj_group_bin_0141 = frame (4k)
frame_gpio_obj_group_bin_0142 = frame (4k)
frame_gpio_obj_group_bin_0143 = frame (4k)
frame_gpio_obj_group_bin_0144 = frame (4k)
frame_gpio_obj_group_bin_0145 = frame (4k)
frame_gpio_obj_group_bin_0146 = frame (4k)
frame_gpio_obj_group_bin_0148 = frame (4k)
frame_gpio_obj_group_bin_0149 = frame (4k)
frame_gpio_obj_group_bin_0150 = frame (4k)
frame_gpio_obj_group_bin_0151 = frame (4k)
frame_gpio_obj_group_bin_0152 = frame (4k)
frame_gpio_obj_group_bin_0153 = frame (4k)
frame_gpio_obj_group_bin_0154 = frame (4k)
frame_gpio_obj_group_bin_0156 = frame (4k)
frame_gpio_obj_group_bin_0157 = frame (4k)
frame_gpio_obj_group_bin_0158 = frame (4k)
frame_gpio_obj_group_bin_0159 = frame (4k)
frame_gpio_obj_group_bin_0160 = frame (4k)
frame_gpio_obj_group_bin_0161 = frame (4k)
frame_gpio_obj_group_bin_0162 = frame (4k)
frame_gpio_obj_group_bin_0163 = frame (4k)
frame_gpio_obj_group_bin_0164 = frame (4k)
frame_gpio_obj_group_bin_0165 = frame (4k)
frame_gpio_obj_group_bin_0166 = frame (4k)
frame_gpio_obj_group_bin_0168 = frame (4k)
frame_gpio_obj_group_bin_0170 = frame (4k)
frame_gpio_obj_group_bin_0171 = frame (4k)
frame_gpio_obj_group_bin_0172 = frame (4k)
frame_gpio_obj_group_bin_0173 = frame (4k)
frame_gpio_obj_group_bin_0174 = frame (4k)
frame_gpio_obj_group_bin_0175 = frame (4k)
frame_gpio_obj_group_bin_0176 = frame (4k)
frame_gpio_obj_group_bin_0177 = frame (4k)
frame_gpio_obj_group_bin_0178 = frame (4k)
frame_gpio_obj_group_bin_0179 = frame (4k)
frame_gpio_obj_group_bin_0180 = frame (4k)
frame_gpio_obj_group_bin_0181 = frame (4k)
frame_gpio_obj_group_bin_0182 = frame (4k)
frame_gpio_obj_group_bin_0183 = frame (4k)
frame_gpio_obj_group_bin_0184 = frame (4k)
frame_gpio_obj_group_bin_0185 = frame (4k)
frame_gpio_obj_group_bin_0186 = frame (4k)
frame_gpio_obj_group_bin_0188 = frame (4k)
frame_gpio_obj_group_bin_0189 = frame (4k)
frame_gpio_obj_group_bin_0190 = frame (4k)
frame_gpio_obj_group_bin_0191 = frame (4k)
frame_gpio_obj_group_bin_0192 = frame (4k)
frame_gpio_obj_group_bin_0193 = frame (4k)
frame_gpio_obj_group_bin_0194 = frame (4k)
frame_gpio_obj_group_bin_0195 = frame (4k)
frame_gpio_obj_group_bin_0196 = frame (4k)
frame_gpio_obj_group_bin_0197 = frame (4k)
frame_gpio_obj_group_bin_0198 = frame (4k)
frame_gpio_obj_group_bin_0199 = frame (4k)
frame_gpio_obj_group_bin_0201 = frame (4k)
frame_gpio_obj_group_bin_0202 = frame (4k)
frame_gpio_obj_group_bin_0203 = frame (4k)
frame_gpio_obj_group_bin_0204 = frame (4k)
frame_gpio_obj_group_bin_0205 = frame (4k)
frame_gpio_obj_group_bin_0206 = frame (4k)
frame_gpio_obj_group_bin_0207 = frame (4k)
frame_gpio_obj_group_bin_0209 = frame (4k)
frame_gpio_obj_group_bin_0211 = frame (4k)
frame_gpio_obj_group_bin_0212 = frame (4k)
frame_gpio_obj_group_bin_0213 = frame (4k)
frame_gpio_obj_group_bin_0214 = frame (4k)
frame_gpio_obj_group_bin_0215 = frame (4k)
frame_gpio_obj_group_bin_0216 = frame (4k)
frame_gpio_obj_group_bin_0217 = frame (4k)
frame_gpio_obj_group_bin_0218 = frame (4k)
frame_gpio_obj_group_bin_0219 = frame (4k)
frame_gpio_obj_group_bin_0220 = frame (4k)
frame_gpio_obj_group_bin_0221 = frame (4k)
frame_gpio_obj_group_bin_0222 = frame (4k)
frame_gpio_obj_group_bin_0223 = frame (4k, paddr: 0x14000000)
frame_gpio_obj_group_bin_0224 = frame (4k)
frame_gpio_obj_group_bin_0225 = frame (4k)
frame_gpio_obj_group_bin_0226 = frame (4k)
frame_gpio_obj_group_bin_0227 = frame (4k)
frame_gpio_obj_group_bin_0228 = frame (4k)
frame_gpio_obj_group_bin_0230 = frame (4k)
frame_gpio_obj_group_bin_0231 = frame (4k)
frame_gpio_obj_group_bin_0232 = frame (4k, paddr: 0x10020000)
frame_gpio_obj_group_bin_0233 = frame (4k)
frame_gpio_obj_group_bin_0234 = frame (4k)
frame_gpio_obj_group_bin_0235 = frame (4k)
frame_gpio_obj_group_bin_0236 = frame (4k)
frame_gpio_obj_group_bin_0237 = frame (4k)
frame_gpio_obj_group_bin_0238 = frame (4k)
frame_gpio_obj_group_bin_0239 = frame (4k)
frame_gpio_obj_group_bin_0240 = frame (4k)
frame_gpio_obj_group_bin_0242 = frame (4k)
frame_gpio_obj_group_bin_0243 = frame (4k)
frame_gpio_obj_group_bin_0244 = frame (4k)
frame_gpio_obj_group_bin_0245 = frame (4k)
frame_gpio_obj_group_bin_0246 = frame (4k)
frame_gpio_obj_group_bin_0247 = frame (4k)
frame_gpio_obj_group_bin_0248 = frame (4k)
frame_gpio_obj_group_bin_0250 = frame (4k)
frame_gpio_obj_group_bin_0252 = frame (4k)
frame_gpio_obj_group_bin_0253 = frame (4k)
frame_gpio_obj_group_bin_0254 = frame (4k)
frame_gpio_obj_group_bin_0255 = frame (4k)
frame_gpio_obj_group_bin_0256 = frame (4k)
frame_gpio_obj_group_bin_0257 = frame (4k)
frame_gpio_obj_group_bin_0258 = frame (4k)
frame_gpio_obj_group_bin_0259 = frame (4k)
frame_gpio_obj_group_bin_0260 = frame (4k)
frame_gpio_obj_group_bin_0261 = frame (4k)
frame_gpio_obj_group_bin_0262 = frame (4k)
frame_gpio_obj_group_bin_0263 = frame (4k)
frame_gpio_obj_group_bin_0264 = frame (4k)
frame_gpio_obj_group_bin_0265 = frame (4k)
frame_gpio_obj_group_bin_0266 = frame (4k)
frame_gpio_obj_group_bin_0267 = frame (4k)
frame_gpio_obj_group_bin_0269 = frame (4k)
frame_gpio_obj_group_bin_0270 = frame (4k)
frame_gpio_obj_group_bin_0271 = frame (4k)
frame_gpio_obj_group_bin_0272 = frame (4k)
frame_gpio_obj_group_bin_0273 = frame (4k)
frame_gpio_obj_group_bin_0274 = frame (4k)
frame_gpio_obj_group_bin_0275 = frame (4k)
frame_gpio_obj_group_bin_0276 = frame (4k)
frame_gpio_obj_group_bin_0277 = frame (4k)
frame_gpio_obj_group_bin_0278 = frame (4k)
frame_gpio_obj_group_bin_0280 = frame (4k)
frame_gpio_obj_group_bin_0281 = frame (4k)
frame_gpio_obj_group_bin_0282 = frame (4k)
frame_gpio_obj_group_bin_0283 = frame (4k)
frame_gpio_obj_group_bin_0285 = frame (4k)
frame_gpio_obj_group_bin_0286 = frame (4k)
frame_gpio_obj_group_bin_0288 = frame (4k)
frame_gpio_obj_group_bin_0289 = frame (4k)
frame_gpio_obj_group_bin_0290 = frame (4k)
frame_gpio_obj_group_bin_0291 = frame (4k)
frame_gpio_obj_group_bin_0292 = frame (4k)
frame_gpio_obj_group_bin_0293 = frame (4k)
frame_gpio_obj_group_bin_0294 = frame (4k)
frame_gpio_obj_group_bin_0295 = frame (4k)
frame_gpio_obj_group_bin_0296 = frame (4k)
frame_gpio_obj_group_bin_0297 = frame (4k)
frame_gpio_obj_group_bin_0298 = frame (4k)
frame_gpio_obj_group_bin_0299 = frame (4k)
frame_gpio_obj_group_bin_0300 = frame (4k)
frame_gpio_obj_group_bin_0301 = frame (4k)
frame_gpio_obj_group_bin_0302 = frame (4k)
frame_gpio_obj_group_bin_0303 = frame (4k)
frame_gpio_obj_group_bin_0304 = frame (4k)
frame_gpio_obj_group_bin_0305 = frame (4k)
frame_gpio_obj_group_bin_0306 = frame (4k)
frame_gpio_obj_group_bin_0307 = frame (4k)
frame_gpio_obj_group_bin_0308 = frame (4k)
frame_gpio_obj_group_bin_0309 = frame (4k)
frame_gpio_obj_group_bin_0310 = frame (4k)
frame_gpio_obj_group_bin_0311 = frame (4k)
frame_gpio_obj_group_bin_0312 = frame (4k)
frame_gpio_obj_group_bin_0313 = frame (4k)
frame_gpio_obj_group_bin_0314 = frame (4k)
frame_gpio_obj_group_bin_0315 = frame (4k)
frame_gpio_obj_group_bin_0316 = frame (4k)
frame_gpio_obj_group_bin_0317 = frame (4k)
frame_gpio_obj_group_bin_0318 = frame (4k)
frame_gpio_obj_group_bin_0319 = frame (4k)
frame_gpio_obj_group_bin_0321 = frame (4k)
frame_gpio_obj_group_bin_0322 = frame (4k)
frame_gpio_obj_group_bin_0323 = frame (4k)
frame_gpio_obj_group_bin_0324 = frame (4k)
frame_gpio_obj_group_bin_0325 = frame (4k)
frame_gpio_obj_group_bin_0326 = frame (4k)
frame_gpio_obj_group_bin_0327 = frame (4k)
frame_gpio_obj_group_bin_0329 = frame (4k)
frame_gpio_obj_group_bin_0330 = frame (4k)
frame_gpio_obj_group_bin_0331 = frame (4k)
frame_gpio_obj_group_bin_0332 = frame (4k)
frame_gpio_obj_group_bin_0333 = frame (4k)
frame_gpio_obj_group_bin_0334 = frame (4k)
frame_gpio_obj_group_bin_0335 = frame (4k)
frame_gpio_obj_group_bin_0336 = frame (4k)
frame_gpio_obj_group_bin_0337 = frame (4k)
frame_gpio_obj_group_bin_0338 = frame (4k)
frame_gpio_obj_group_bin_0339 = frame (4k)
frame_gpio_obj_group_bin_0340 = frame (4k)
frame_gpio_obj_group_bin_0341 = frame (4k)
frame_gpio_obj_group_bin_0342 = frame (4k)
frame_gpio_obj_group_bin_0343 = frame (4k)
frame_gpio_obj_group_bin_0344 = frame (4k)
frame_gpio_obj_group_bin_0345 = frame (4k)
frame_gpio_obj_group_bin_0346 = frame (4k)
frame_gpio_obj_group_bin_0347 = frame (4k)
frame_gpio_obj_group_bin_0348 = frame (4k)
frame_gpio_obj_group_bin_0349 = frame (4k)
frame_gpio_obj_group_bin_0350 = frame (4k)
frame_gpio_obj_group_bin_0351 = frame (4k)
frame_gpio_obj_group_bin_0352 = frame (4k)
frame_gpio_obj_group_bin_0353 = frame (4k)
frame_gpio_obj_group_bin_0354 = frame (4k)
frame_gpio_obj_group_bin_0355 = frame (4k)
frame_pilot_obj_group_bin_0000 = frame (4k)
frame_pilot_obj_group_bin_0001 = frame (4k)
frame_pilot_obj_group_bin_0002 = frame (4k)
frame_pilot_obj_group_bin_0003 = frame (4k)
frame_pilot_obj_group_bin_0004 = frame (4k)
frame_pilot_obj_group_bin_0005 = frame (4k)
frame_pilot_obj_group_bin_0006 = frame (4k)
frame_pilot_obj_group_bin_0007 = frame (4k)
frame_pilot_obj_group_bin_0008 = frame (4k)
frame_pilot_obj_group_bin_0009 = frame (4k)
frame_pilot_obj_group_bin_0010 = frame (4k)
frame_pilot_obj_group_bin_0011 = frame (4k)
frame_pilot_obj_group_bin_0012 = frame (4k)
frame_pilot_obj_group_bin_0013 = frame (4k)
frame_pilot_obj_group_bin_0014 = frame (4k)
frame_pilot_obj_group_bin_0015 = frame (4k)
frame_pilot_obj_group_bin_0016 = frame (4k)
frame_pilot_obj_group_bin_0017 = frame (4k)
frame_pilot_obj_group_bin_0018 = frame (4k)
frame_pilot_obj_group_bin_0019 = frame (4k)
frame_pilot_obj_group_bin_0020 = frame (4k)
frame_pilot_obj_group_bin_0021 = frame (4k)
frame_pilot_obj_group_bin_0022 = frame (4k)
frame_pilot_obj_group_bin_0023 = frame (4k)
frame_pilot_obj_group_bin_0024 = frame (4k)
frame_pilot_obj_group_bin_0025 = frame (4k)
frame_pilot_obj_group_bin_0026 = frame (4k)
frame_pilot_obj_group_bin_0027 = frame (4k)
frame_pilot_obj_group_bin_0029 = frame (4k)
frame_pilot_obj_group_bin_0030 = frame (4k)
frame_pilot_obj_group_bin_0031 = frame (4k)
frame_pilot_obj_group_bin_0032 = frame (4k)
frame_pilot_obj_group_bin_0033 = frame (4k)
frame_pilot_obj_group_bin_0034 = frame (4k)
frame_pilot_obj_group_bin_0035 = frame (4k)
frame_pilot_obj_group_bin_0036 = frame (4k)
frame_pilot_obj_group_bin_0037 = frame (4k)
frame_pilot_obj_group_bin_0038 = frame (4k)
frame_pilot_obj_group_bin_0039 = frame (4k)
frame_pilot_obj_group_bin_0040 = frame (4k)
frame_pilot_obj_group_bin_0042 = frame (4k)
frame_pilot_obj_group_bin_0043 = frame (4k)
frame_pilot_obj_group_bin_0044 = frame (4k)
frame_pilot_obj_group_bin_0045 = frame (4k)
frame_pilot_obj_group_bin_0046 = frame (4k)
frame_pilot_obj_group_bin_0047 = frame (4k)
frame_pilot_obj_group_bin_0048 = frame (4k)
frame_pilot_obj_group_bin_0049 = frame (4k)
frame_pilot_obj_group_bin_0050 = frame (4k)
frame_pilot_obj_group_bin_0051 = frame (4k)
frame_pilot_obj_group_bin_0052 = frame (4k)
frame_pilot_obj_group_bin_0053 = frame (4k)
frame_pilot_obj_group_bin_0054 = frame (4k)
frame_pilot_obj_group_bin_0055 = frame (4k)
frame_pilot_obj_group_bin_0056 = frame (4k)
frame_pilot_obj_group_bin_0057 = frame (4k)
frame_pilot_obj_group_bin_0058 = frame (4k)
frame_pilot_obj_group_bin_0059 = frame (4k)
frame_pilot_obj_group_bin_0060 = frame (4k)
frame_pilot_obj_group_bin_0061 = frame (4k)
frame_pilot_obj_group_bin_0062 = frame (4k)
frame_pilot_obj_group_bin_0064 = frame (4k)
frame_pilot_obj_group_bin_0065 = frame (4k)
frame_pilot_obj_group_bin_0066 = frame (4k)
frame_pilot_obj_group_bin_0067 = frame (4k)
frame_pilot_obj_group_bin_0068 = frame (4k)
frame_pilot_obj_group_bin_0069 = frame (4k)
frame_pilot_obj_group_bin_0070 = frame (4k)
frame_pilot_obj_group_bin_0071 = frame (4k)
frame_pilot_obj_group_bin_0072 = frame (4k)
frame_pilot_obj_group_bin_0073 = frame (4k)
frame_pilot_obj_group_bin_0074 = frame (4k)
frame_pilot_obj_group_bin_0075 = frame (4k)
frame_pilot_obj_group_bin_0076 = frame (4k)
frame_pilot_obj_group_bin_0077 = frame (4k)
frame_pilot_obj_group_bin_0078 = frame (4k)
frame_pilot_obj_group_bin_0079 = frame (4k)
frame_pilot_obj_group_bin_0080 = frame (4k)
frame_pilot_obj_group_bin_0081 = frame (4k)
frame_pilot_obj_group_bin_0082 = frame (4k)
frame_pilot_obj_group_bin_0083 = frame (4k)
frame_pilot_obj_group_bin_0084 = frame (4k)
frame_pilot_obj_group_bin_0085 = frame (4k)
frame_pilot_obj_group_bin_0086 = frame (4k)
frame_pilot_obj_group_bin_0087 = frame (4k)
frame_pilot_obj_group_bin_0088 = frame (4k)
frame_pilot_obj_group_bin_0089 = frame (4k)
frame_pilot_obj_group_bin_0090 = frame (4k)
frame_pilot_obj_group_bin_0091 = frame (4k)
frame_pilot_obj_group_bin_0092 = frame (4k)
frame_pilot_obj_group_bin_0093 = frame (4k)
frame_pilot_obj_group_bin_0094 = frame (4k)
frame_pilot_obj_group_bin_0095 = frame (4k)
frame_pilot_obj_group_bin_0096 = frame (4k)
frame_pilot_obj_group_bin_0097 = frame (4k)
frame_pilot_obj_group_bin_0098 = frame (4k)
frame_pilot_obj_group_bin_0099 = frame (4k)
frame_pilot_obj_group_bin_0100 = frame (4k)
frame_pilot_obj_group_bin_0101 = frame (4k)
frame_pilot_obj_group_bin_0102 = frame (4k)
frame_pilot_obj_group_bin_0103 = frame (4k)
frame_pilot_obj_group_bin_0104 = frame (4k)
frame_pilot_obj_group_bin_0105 = frame (4k)
frame_pilot_obj_group_bin_0106 = frame (4k)
frame_pilot_obj_group_bin_0107 = frame (4k)
frame_pilot_obj_group_bin_0108 = frame (4k)
frame_pilot_obj_group_bin_0109 = frame (4k)
frame_pilot_obj_group_bin_0110 = frame (4k)
frame_pilot_obj_group_bin_0112 = frame (4k)
frame_pilot_obj_group_bin_0113 = frame (4k)
frame_pilot_obj_group_bin_0114 = frame (4k)
frame_pilot_obj_group_bin_0115 = frame (4k)
frame_pilot_obj_group_bin_0116 = frame (4k)
frame_pilot_obj_group_bin_0117 = frame (4k)
frame_pilot_obj_group_bin_0119 = frame (4k)
frame_pilot_obj_group_bin_0120 = frame (4k)
frame_pilot_obj_group_bin_0121 = frame (4k)
frame_pilot_obj_group_bin_0122 = frame (4k)
frame_pilot_obj_group_bin_0123 = frame (4k)
frame_pilot_obj_group_bin_0124 = frame (4k)
frame_pilot_obj_group_bin_0125 = frame (4k)
frame_pilot_obj_group_bin_0126 = frame (4k)
frame_pilot_obj_group_bin_0127 = frame (4k)
frame_pilot_obj_group_bin_0128 = frame (4k)
frame_pilot_obj_group_bin_0129 = frame (4k)
frame_pilot_obj_group_bin_0130 = frame (4k)
frame_pilot_obj_group_bin_0132 = frame (4k)
frame_pilot_obj_group_bin_0133 = frame (4k)
frame_pilot_obj_group_bin_0134 = frame (4k)
frame_pilot_obj_group_bin_0135 = frame (4k)
frame_pilot_obj_group_bin_0136 = frame (4k)
frame_pilot_obj_group_bin_0137 = frame (4k)
frame_pilot_obj_group_bin_0138 = frame (4k)
frame_pilot_obj_group_bin_0139 = frame (4k)
frame_pilot_obj_group_bin_0140 = frame (4k)
frame_pilot_obj_group_bin_0141 = frame (4k)
frame_pilot_obj_group_bin_0143 = frame (4k)
frame_pilot_obj_group_bin_0144 = frame (4k)
frame_pilot_obj_group_bin_0145 = frame (4k)
frame_pilot_obj_group_bin_0146 = frame (4k)
frame_pilot_obj_group_bin_0147 = frame (4k)
frame_pilot_obj_group_bin_0148 = frame (4k)
frame_pilot_obj_group_bin_0149 = frame (4k)
frame_pilot_obj_group_bin_0150 = frame (4k)
frame_pilot_obj_group_bin_0151 = frame (4k)
frame_pilot_obj_group_bin_0152 = frame (4k)
frame_pilot_obj_group_bin_0153 = frame (4k)
frame_pilot_obj_group_bin_0154 = frame (4k)
frame_pilot_obj_group_bin_0155 = frame (4k)
frame_pilot_obj_group_bin_0156 = frame (4k)
frame_pilot_obj_group_bin_0157 = frame (4k)
frame_pilot_obj_group_bin_0158 = frame (4k)
frame_pilot_obj_group_bin_0159 = frame (4k)
frame_pilot_obj_group_bin_0160 = frame (4k)
frame_pilot_obj_group_bin_0161 = frame (4k)
frame_pilot_obj_group_bin_0162 = frame (4k)
frame_pilot_obj_group_bin_0163 = frame (4k)
frame_pilot_obj_group_bin_0164 = frame (4k)
frame_pilot_obj_group_bin_0165 = frame (4k)
frame_pilot_obj_group_bin_0166 = frame (4k)
frame_pilot_obj_group_bin_0167 = frame (4k)
frame_pilot_obj_group_bin_0168 = frame (4k)
frame_pilot_obj_group_bin_0169 = frame (4k)
frame_pilot_obj_group_bin_0170 = frame (4k)
frame_pilot_obj_group_bin_0171 = frame (4k)
frame_pilot_obj_group_bin_0172 = frame (4k)
frame_pilot_obj_group_bin_0173 = frame (4k)
frame_pilot_obj_group_bin_0174 = frame (4k)
frame_pilot_obj_group_bin_0175 = frame (4k)
frame_pilot_obj_group_bin_0176 = frame (4k)
frame_pilot_obj_group_bin_0177 = frame (4k)
frame_pilot_obj_group_bin_0178 = frame (4k)
frame_pilot_obj_group_bin_0179 = frame (4k)
frame_pilot_obj_group_bin_0180 = frame (4k)
frame_pilot_obj_group_bin_0181 = frame (4k)
frame_pilot_obj_group_bin_0182 = frame (4k)
frame_pilot_obj_group_bin_0183 = frame (4k)
frame_pilot_obj_group_bin_0184 = frame (4k)
frame_pilot_obj_group_bin_0185 = frame (4k)
frame_pilot_obj_group_bin_0186 = frame (4k)
frame_pilot_obj_group_bin_0187 = frame (4k)
frame_pilot_obj_group_bin_0189 = frame (4k)
frame_pilot_obj_group_bin_0190 = frame (4k)
frame_pilot_obj_group_bin_0191 = frame (4k)
frame_pilot_obj_group_bin_0192 = frame (4k)
frame_pilot_obj_group_bin_0193 = frame (4k)
frame_pilot_obj_group_bin_0194 = frame (4k)
frame_pilot_obj_group_bin_0195 = frame (4k)
frame_pilot_obj_group_bin_0196 = frame (4k)
frame_pilot_obj_group_bin_0197 = frame (4k)
frame_pilot_obj_group_bin_0198 = frame (4k)
frame_pilot_obj_group_bin_0199 = frame (4k)
frame_pilot_obj_group_bin_0200 = frame (4k)
frame_pilot_obj_group_bin_0201 = frame (4k)
frame_pilot_obj_group_bin_0202 = frame (4k)
frame_pilot_obj_group_bin_0203 = frame (4k)
frame_pilot_obj_group_bin_0204 = frame (4k)
frame_pilot_obj_group_bin_0205 = frame (4k)
frame_pilot_obj_group_bin_0207 = frame (4k)
frame_pilot_obj_group_bin_0208 = frame (4k)
frame_pilot_obj_group_bin_0209 = frame (4k)
frame_pilot_obj_group_bin_0210 = frame (4k)
frame_pilot_obj_group_bin_0211 = frame (4k)
frame_pilot_obj_group_bin_0212 = frame (4k)
frame_pilot_obj_group_bin_0213 = frame (4k)
frame_pilot_obj_group_bin_0214 = frame (4k)
frame_pilot_obj_group_bin_0215 = frame (4k)
frame_pilot_obj_group_bin_0216 = frame (4k)
frame_pilot_obj_group_bin_0217 = frame (4k)
frame_pilot_obj_group_bin_0218 = frame (4k)
frame_pilot_obj_group_bin_0219 = frame (4k)
frame_pilot_obj_group_bin_0220 = frame (4k)
frame_pilot_obj_group_bin_0221 = frame (4k)
frame_pilot_obj_group_bin_0222 = frame (4k)
frame_pilot_obj_group_bin_0223 = frame (4k)
frame_pilot_obj_group_bin_0224 = frame (4k)
frame_pilot_obj_group_bin_0225 = frame (4k)
frame_pilot_obj_group_bin_0226 = frame (4k)
frame_pilot_obj_group_bin_0227 = frame (4k)
frame_pilot_obj_group_bin_0228 = frame (4k)
frame_pilot_obj_group_bin_0229 = frame (4k)
frame_pilot_obj_group_bin_0230 = frame (4k)
frame_pilot_obj_group_bin_0231 = frame (4k)
frame_pilot_obj_group_bin_0232 = frame (4k)
frame_pilot_obj_group_bin_0233 = frame (4k)
frame_pilot_obj_group_bin_0234 = frame (4k)
frame_pilot_obj_group_bin_0235 = frame (4k)
frame_pilot_obj_group_bin_0236 = frame (4k)
frame_pilot_obj_group_bin_0237 = frame (4k)
frame_pilot_obj_group_bin_0238 = frame (4k)
frame_pilot_obj_group_bin_0239 = frame (4k)
frame_pilot_obj_group_bin_0240 = frame (4k)
frame_pilot_obj_group_bin_0242 = frame (4k)
frame_pilot_obj_group_bin_0243 = frame (4k)
frame_pilot_obj_group_bin_0244 = frame (4k)
frame_pilot_obj_group_bin_0245 = frame (4k)
frame_pilot_obj_group_bin_0246 = frame (4k)
frame_pilot_obj_group_bin_0247 = frame (4k)
frame_pilot_obj_group_bin_0248 = frame (4k)
frame_pilot_obj_group_bin_0249 = frame (4k)
frame_pilot_obj_group_bin_0250 = frame (4k)
frame_pilot_obj_group_bin_0251 = frame (4k)
frame_pilot_obj_group_bin_0252 = frame (4k)
frame_pilot_obj_group_bin_0253 = frame (4k)
frame_pilot_obj_group_bin_0254 = frame (4k)
frame_pilot_obj_group_bin_0255 = frame (4k)
frame_pilot_obj_group_bin_0256 = frame (4k)
frame_pilot_obj_group_bin_0257 = frame (4k)
frame_pilot_obj_group_bin_0258 = frame (4k)
frame_pilot_obj_group_bin_0259 = frame (4k)
frame_pilot_obj_group_bin_0260 = frame (4k)
frame_pilot_obj_group_bin_0261 = frame (4k)
frame_pilot_obj_group_bin_0262 = frame (4k)
frame_pilot_obj_group_bin_0263 = frame (4k)
frame_pilot_obj_group_bin_0264 = frame (4k)
frame_pilot_obj_group_bin_0265 = frame (4k)
frame_pilot_obj_group_bin_0266 = frame (4k)
frame_pilot_obj_group_bin_0267 = frame (4k)
frame_pilot_obj_group_bin_0268 = frame (4k)
frame_pilot_obj_group_bin_0269 = frame (4k)
frame_pilot_obj_group_bin_0270 = frame (4k)
frame_pilot_obj_group_bin_0272 = frame (4k)
frame_pilot_obj_group_bin_0273 = frame (4k)
frame_pilot_obj_group_bin_0274 = frame (4k)
frame_pilot_obj_group_bin_0275 = frame (4k)
frame_pilot_obj_group_bin_0276 = frame (4k)
frame_pilot_obj_group_bin_0277 = frame (4k)
frame_pilot_obj_group_bin_0278 = frame (4k)
frame_pilot_obj_group_bin_0279 = frame (4k)
frame_pilot_obj_group_bin_0280 = frame (4k)
frame_pilot_obj_group_bin_0281 = frame (4k)
frame_pilot_obj_group_bin_0282 = frame (4k)
frame_pilot_obj_group_bin_0283 = frame (4k)
frame_pilot_obj_group_bin_0284 = frame (4k)
frame_pilot_obj_group_bin_0285 = frame (4k)
frame_pilot_obj_group_bin_0286 = frame (4k)
frame_pilot_obj_group_bin_0288 = frame (4k)
frame_pilot_obj_group_bin_0290 = frame (4k)
frame_pilot_obj_group_bin_0291 = frame (4k)
frame_pilot_obj_group_bin_0292 = frame (4k)
frame_pilot_obj_group_bin_0293 = frame (4k)
frame_pilot_obj_group_bin_0294 = frame (4k)
frame_pilot_obj_group_bin_0295 = frame (4k)
frame_pilot_obj_group_bin_0296 = frame (4k)
frame_pilot_obj_group_bin_0297 = frame (4k)
frame_pilot_obj_group_bin_0298 = frame (4k)
frame_pilot_obj_group_bin_0299 = frame (4k)
frame_pilot_obj_group_bin_0300 = frame (4k)
frame_pilot_obj_group_bin_0301 = frame (4k)
frame_pilot_obj_group_bin_0302 = frame (4k)
frame_pilot_obj_group_bin_0303 = frame (4k)
frame_pilot_obj_group_bin_0304 = frame (4k)
frame_pilot_obj_group_bin_0305 = frame (4k)
frame_pilot_obj_group_bin_0306 = frame (4k)
frame_pilot_obj_group_bin_0307 = frame (4k)
frame_pilot_obj_group_bin_0308 = frame (4k)
frame_pilot_obj_group_bin_0309 = frame (4k)
frame_pilot_obj_group_bin_0310 = frame (4k)
frame_pilot_obj_group_bin_0311 = frame (4k)
frame_pilot_obj_group_bin_0312 = frame (4k)
frame_pilot_obj_group_bin_0313 = frame (4k)
frame_pilot_obj_group_bin_0314 = frame (4k)
frame_pilot_obj_group_bin_0315 = frame (4k)
frame_pwm_obj_group_bin_0000 = frame (4k)
frame_pwm_obj_group_bin_0001 = frame (4k)
frame_pwm_obj_group_bin_0002 = frame (4k)
frame_pwm_obj_group_bin_0003 = frame (4k)
frame_pwm_obj_group_bin_0004 = frame (4k)
frame_pwm_obj_group_bin_0005 = frame (4k)
frame_pwm_obj_group_bin_0006 = frame (4k)
frame_pwm_obj_group_bin_0007 = frame (4k)
frame_pwm_obj_group_bin_0008 = frame (4k)
frame_pwm_obj_group_bin_0010 = frame (4k)
frame_pwm_obj_group_bin_0011 = frame (4k)
frame_pwm_obj_group_bin_0012 = frame (4k)
frame_pwm_obj_group_bin_0013 = frame (4k)
frame_pwm_obj_group_bin_0014 = frame (4k)
frame_pwm_obj_group_bin_0015 = frame (4k)
frame_pwm_obj_group_bin_0016 = frame (4k)
frame_pwm_obj_group_bin_0017 = frame (4k)
frame_pwm_obj_group_bin_0018 = frame (4k)
frame_pwm_obj_group_bin_0019 = frame (4k)
frame_pwm_obj_group_bin_0020 = frame (4k)
frame_pwm_obj_group_bin_0021 = frame (4k)
frame_pwm_obj_group_bin_0022 = frame (4k)
frame_pwm_obj_group_bin_0023 = frame (4k)
frame_pwm_obj_group_bin_0024 = frame (4k)
frame_pwm_obj_group_bin_0025 = frame (4k)
frame_pwm_obj_group_bin_0026 = frame (4k)
frame_pwm_obj_group_bin_0028 = frame (4k)
frame_pwm_obj_group_bin_0029 = frame (4k)
frame_pwm_obj_group_bin_0030 = frame (4k)
frame_pwm_obj_group_bin_0031 = frame (4k)
frame_pwm_obj_group_bin_0032 = frame (4k)
frame_pwm_obj_group_bin_0033 = frame (4k)
frame_pwm_obj_group_bin_0034 = frame (4k)
frame_pwm_obj_group_bin_0035 = frame (4k)
frame_pwm_obj_group_bin_0036 = frame (4k)
frame_pwm_obj_group_bin_0037 = frame (4k)
frame_pwm_obj_group_bin_0038 = frame (4k)
frame_pwm_obj_group_bin_0039 = frame (4k)
frame_pwm_obj_group_bin_0040 = frame (4k)
frame_pwm_obj_group_bin_0041 = frame (4k)
frame_pwm_obj_group_bin_0042 = frame (4k)
frame_pwm_obj_group_bin_0043 = frame (4k)
frame_pwm_obj_group_bin_0044 = frame (4k)
frame_pwm_obj_group_bin_0045 = frame (4k)
frame_pwm_obj_group_bin_0046 = frame (4k)
frame_pwm_obj_group_bin_0047 = frame (4k)
frame_pwm_obj_group_bin_0048 = frame (4k)
frame_pwm_obj_group_bin_0049 = frame (4k)
frame_pwm_obj_group_bin_0050 = frame (4k)
frame_pwm_obj_group_bin_0051 = frame (4k)
frame_pwm_obj_group_bin_0052 = frame (4k)
frame_pwm_obj_group_bin_0053 = frame (4k)
frame_pwm_obj_group_bin_0054 = frame (4k)
frame_pwm_obj_group_bin_0055 = frame (4k)
frame_pwm_obj_group_bin_0056 = frame (4k)
frame_pwm_obj_group_bin_0057 = frame (4k)
frame_pwm_obj_group_bin_0058 = frame (4k)
frame_pwm_obj_group_bin_0059 = frame (4k)
frame_pwm_obj_group_bin_0060 = frame (4k)
frame_pwm_obj_group_bin_0061 = frame (4k)
frame_pwm_obj_group_bin_0062 = frame (4k)
frame_pwm_obj_group_bin_0063 = frame (4k)
frame_pwm_obj_group_bin_0064 = frame (4k)
frame_pwm_obj_group_bin_0065 = frame (4k)
frame_pwm_obj_group_bin_0067 = frame (4k)
frame_pwm_obj_group_bin_0068 = frame (4k)
frame_pwm_obj_group_bin_0069 = frame (4k)
frame_pwm_obj_group_bin_0070 = frame (4k)
frame_pwm_obj_group_bin_0071 = frame (4k)
frame_pwm_obj_group_bin_0072 = frame (4k)
frame_pwm_obj_group_bin_0073 = frame (4k)
frame_pwm_obj_group_bin_0074 = frame (4k)
frame_pwm_obj_group_bin_0075 = frame (4k)
frame_pwm_obj_group_bin_0076 = frame (4k)
frame_pwm_obj_group_bin_0077 = frame (4k)
frame_pwm_obj_group_bin_0078 = frame (4k)
frame_pwm_obj_group_bin_0079 = frame (4k)
frame_pwm_obj_group_bin_0080 = frame (4k)
frame_pwm_obj_group_bin_0081 = frame (4k)
frame_pwm_obj_group_bin_0082 = frame (4k)
frame_pwm_obj_group_bin_0083 = frame (4k)
frame_pwm_obj_group_bin_0084 = frame (4k)
frame_pwm_obj_group_bin_0085 = frame (4k)
frame_pwm_obj_group_bin_0086 = frame (4k)
frame_pwm_obj_group_bin_0087 = frame (4k)
frame_pwm_obj_group_bin_0088 = frame (4k)
frame_pwm_obj_group_bin_0089 = frame (4k)
frame_pwm_obj_group_bin_0090 = frame (4k)
frame_pwm_obj_group_bin_0092 = frame (4k)
frame_pwm_obj_group_bin_0093 = frame (4k)
frame_pwm_obj_group_bin_0094 = frame (4k)
frame_pwm_obj_group_bin_0095 = frame (4k)
frame_pwm_obj_group_bin_0096 = frame (4k)
frame_pwm_obj_group_bin_0097 = frame (4k)
frame_pwm_obj_group_bin_0098 = frame (4k)
frame_pwm_obj_group_bin_0099 = frame (4k)
frame_pwm_obj_group_bin_0100 = frame (4k)
frame_pwm_obj_group_bin_0102 = frame (4k)
frame_pwm_obj_group_bin_0103 = frame (4k)
frame_pwm_obj_group_bin_0104 = frame (4k)
frame_pwm_obj_group_bin_0105 = frame (4k)
frame_pwm_obj_group_bin_0106 = frame (4k)
frame_pwm_obj_group_bin_0107 = frame (4k)
frame_pwm_obj_group_bin_0109 = frame (4k)
frame_pwm_obj_group_bin_0110 = frame (4k)
frame_pwm_obj_group_bin_0111 = frame (4k)
frame_pwm_obj_group_bin_0112 = frame (4k)
frame_pwm_obj_group_bin_0114 = frame (4k)
frame_pwm_obj_group_bin_0115 = frame (4k)
frame_pwm_obj_group_bin_0116 = frame (4k)
frame_pwm_obj_group_bin_0117 = frame (4k)
frame_pwm_obj_group_bin_0118 = frame (4k)
frame_pwm_obj_group_bin_0119 = frame (4k)
frame_pwm_obj_group_bin_0120 = frame (4k)
frame_pwm_obj_group_bin_0121 = frame (4k)
frame_pwm_obj_group_bin_0122 = frame (4k)
frame_pwm_obj_group_bin_0123 = frame (4k)
frame_pwm_obj_group_bin_0124 = frame (4k)
frame_pwm_obj_group_bin_0125 = frame (4k)
frame_pwm_obj_group_bin_0126 = frame (4k)
frame_pwm_obj_group_bin_0127 = frame (4k)
frame_pwm_obj_group_bin_0128 = frame (4k)
frame_pwm_obj_group_bin_0129 = frame (4k)
frame_pwm_obj_group_bin_0130 = frame (4k)
frame_pwm_obj_group_bin_0131 = frame (4k)
frame_pwm_obj_group_bin_0132 = frame (4k)
frame_pwm_obj_group_bin_0133 = frame (4k)
frame_pwm_obj_group_bin_0134 = frame (4k)
frame_pwm_obj_group_bin_0135 = frame (4k)
frame_pwm_obj_group_bin_0136 = frame (4k)
frame_pwm_obj_group_bin_0138 = frame (4k)
frame_pwm_obj_group_bin_0139 = frame (4k)
frame_pwm_obj_group_bin_0140 = frame (4k)
frame_pwm_obj_group_bin_0141 = frame (4k)
frame_pwm_obj_group_bin_0142 = frame (4k)
frame_pwm_obj_group_bin_0143 = frame (4k)
frame_pwm_obj_group_bin_0144 = frame (4k)
frame_pwm_obj_group_bin_0145 = frame (4k)
frame_pwm_obj_group_bin_0146 = frame (4k)
frame_pwm_obj_group_bin_0147 = frame (4k)
frame_pwm_obj_group_bin_0148 = frame (4k)
frame_pwm_obj_group_bin_0150 = frame (4k)
frame_pwm_obj_group_bin_0151 = frame (4k)
frame_pwm_obj_group_bin_0152 = frame (4k)
frame_pwm_obj_group_bin_0153 = frame (4k)
frame_pwm_obj_group_bin_0154 = frame (4k)
frame_pwm_obj_group_bin_0156 = frame (4k)
frame_pwm_obj_group_bin_0157 = frame (4k)
frame_pwm_obj_group_bin_0158 = frame (4k)
frame_pwm_obj_group_bin_0159 = frame (4k)
frame_pwm_obj_group_bin_0162 = frame (4k)
frame_pwm_obj_group_bin_0163 = frame (4k)
frame_pwm_obj_group_bin_0164 = frame (4k)
frame_pwm_obj_group_bin_0165 = frame (4k)
frame_pwm_obj_group_bin_0166 = frame (4k)
frame_pwm_obj_group_bin_0167 = frame (4k)
frame_pwm_obj_group_bin_0168 = frame (4k)
frame_pwm_obj_group_bin_0169 = frame (4k)
frame_pwm_obj_group_bin_0170 = frame (4k)
frame_pwm_obj_group_bin_0171 = frame (4k)
frame_pwm_obj_group_bin_0172 = frame (4k)
frame_pwm_obj_group_bin_0173 = frame (4k)
frame_pwm_obj_group_bin_0174 = frame (4k)
frame_pwm_obj_group_bin_0175 = frame (4k)
frame_pwm_obj_group_bin_0176 = frame (4k)
frame_pwm_obj_group_bin_0177 = frame (4k)
frame_pwm_obj_group_bin_0178 = frame (4k)
frame_pwm_obj_group_bin_0179 = frame (4k)
frame_pwm_obj_group_bin_0181 = frame (4k)
frame_pwm_obj_group_bin_0182 = frame (4k)
frame_pwm_obj_group_bin_0183 = frame (4k)
frame_pwm_obj_group_bin_0184 = frame (4k)
frame_pwm_obj_group_bin_0185 = frame (4k)
frame_pwm_obj_group_bin_0186 = frame (4k)
frame_pwm_obj_group_bin_0187 = frame (4k)
frame_pwm_obj_group_bin_0188 = frame (4k)
frame_pwm_obj_group_bin_0189 = frame (4k)
frame_pwm_obj_group_bin_0190 = frame (4k)
frame_pwm_obj_group_bin_0191 = frame (4k)
frame_pwm_obj_group_bin_0192 = frame (4k)
frame_pwm_obj_group_bin_0193 = frame (4k)
frame_pwm_obj_group_bin_0194 = frame (4k)
frame_pwm_obj_group_bin_0195 = frame (4k)
frame_pwm_obj_group_bin_0196 = frame (4k)
frame_pwm_obj_group_bin_0197 = frame (4k)
frame_pwm_obj_group_bin_0198 = frame (4k)
frame_pwm_obj_group_bin_0199 = frame (4k)
frame_pwm_obj_group_bin_0200 = frame (4k)
frame_pwm_obj_group_bin_0201 = frame (4k)
frame_pwm_obj_group_bin_0202 = frame (4k)
frame_pwm_obj_group_bin_0203 = frame (4k)
frame_pwm_obj_group_bin_0204 = frame (4k)
frame_pwm_obj_group_bin_0205 = frame (4k)
frame_pwm_obj_group_bin_0206 = frame (4k)
frame_pwm_obj_group_bin_0207 = frame (4k)
frame_pwm_obj_group_bin_0209 = frame (4k)
frame_pwm_obj_group_bin_0210 = frame (4k)
frame_pwm_obj_group_bin_0213 = frame (4k)
frame_pwm_obj_group_bin_0214 = frame (4k)
frame_pwm_obj_group_bin_0215 = frame (4k)
frame_pwm_obj_group_bin_0216 = frame (4k)
frame_pwm_obj_group_bin_0217 = frame (4k)
frame_pwm_obj_group_bin_0218 = frame (4k)
frame_pwm_obj_group_bin_0219 = frame (4k)
frame_pwm_obj_group_bin_0220 = frame (4k)
frame_pwm_obj_group_bin_0221 = frame (4k)
frame_pwm_obj_group_bin_0222 = frame (4k)
frame_pwm_obj_group_bin_0223 = frame (4k)
frame_pwm_obj_group_bin_0224 = frame (4k)
frame_pwm_obj_group_bin_0225 = frame (4k)
frame_pwm_obj_group_bin_0226 = frame (4k)
frame_pwm_obj_group_bin_0227 = frame (4k)
frame_pwm_obj_group_bin_0228 = frame (4k)
frame_pwm_obj_group_bin_0229 = frame (4k)
frame_pwm_obj_group_bin_0230 = frame (4k)
frame_pwm_obj_group_bin_0231 = frame (4k)
frame_pwm_obj_group_bin_0232 = frame (4k)
frame_pwm_obj_group_bin_0233 = frame (4k)
frame_pwm_obj_group_bin_0235 = frame (4k)
frame_pwm_obj_group_bin_0236 = frame (4k)
frame_pwm_obj_group_bin_0237 = frame (4k)
frame_pwm_obj_group_bin_0238 = frame (4k)
frame_pwm_obj_group_bin_0239 = frame (4k)
frame_pwm_obj_group_bin_0240 = frame (4k)
frame_pwm_obj_group_bin_0241 = frame (4k)
frame_pwm_obj_group_bin_0242 = frame (4k)
frame_pwm_obj_group_bin_0243 = frame (4k)
frame_pwm_obj_group_bin_0244 = frame (4k)
frame_pwm_obj_group_bin_0246 = frame (4k)
frame_pwm_obj_group_bin_0247 = frame (4k)
frame_pwm_obj_group_bin_0248 = frame (4k)
frame_pwm_obj_group_bin_0249 = frame (4k)
frame_pwm_obj_group_bin_0250 = frame (4k)
frame_pwm_obj_group_bin_0252 = frame (4k)
frame_pwm_obj_group_bin_0253 = frame (4k)
frame_pwm_obj_group_bin_0254 = frame (4k)
frame_pwm_obj_group_bin_0255 = frame (4k)
frame_pwm_obj_group_bin_0256 = frame (4k)
frame_pwm_obj_group_bin_0257 = frame (4k)
frame_pwm_obj_group_bin_0258 = frame (4k, paddr: 0x12c60000)
frame_pwm_obj_group_bin_0259 = frame (4k)
frame_pwm_obj_group_bin_0260 = frame (4k)
frame_pwm_obj_group_bin_0261 = frame (4k)
frame_pwm_obj_group_bin_0262 = frame (4k)
frame_pwm_obj_group_bin_0263 = frame (4k)
frame_pwm_obj_group_bin_0265 = frame (4k)
frame_pwm_obj_group_bin_0266 = frame (4k)
frame_pwm_obj_group_bin_0267 = frame (4k)
frame_pwm_obj_group_bin_0268 = frame (4k)
frame_pwm_obj_group_bin_0269 = frame (4k)
frame_pwm_obj_group_bin_0270 = frame (4k)
frame_pwm_obj_group_bin_0271 = frame (4k)
frame_pwm_obj_group_bin_0273 = frame (4k)
frame_pwm_obj_group_bin_0275 = frame (4k)
frame_pwm_obj_group_bin_0277 = frame (4k)
frame_pwm_obj_group_bin_0278 = frame (4k)
frame_pwm_obj_group_bin_0279 = frame (4k)
frame_pwm_obj_group_bin_0280 = frame (4k)
frame_pwm_obj_group_bin_0281 = frame (4k)
frame_pwm_obj_group_bin_0282 = frame (4k)
frame_pwm_obj_group_bin_0283 = frame (4k)
frame_pwm_obj_group_bin_0284 = frame (4k)
frame_pwm_obj_group_bin_0285 = frame (4k)
frame_pwm_obj_group_bin_0286 = frame (4k)
frame_pwm_obj_group_bin_0287 = frame (4k)
frame_pwm_obj_group_bin_0288 = frame (4k)
frame_pwm_obj_group_bin_0289 = frame (4k)
frame_pwm_obj_group_bin_0290 = frame (4k)
frame_pwm_obj_group_bin_0291 = frame (4k)
frame_pwm_obj_group_bin_0292 = frame (4k)
frame_pwm_obj_group_bin_0293 = frame (4k)
frame_pwm_obj_group_bin_0294 = frame (4k)
frame_pwm_obj_group_bin_0295 = frame (4k)
frame_pwm_obj_group_bin_0296 = frame (4k)
frame_pwm_obj_group_bin_0297 = frame (4k)
frame_pwm_obj_group_bin_0298 = frame (4k)
frame_pwm_obj_group_bin_0299 = frame (4k)
frame_pwm_obj_group_bin_0300 = frame (4k)
frame_pwm_obj_group_bin_0301 = frame (4k)
frame_pwm_obj_group_bin_0302 = frame (4k)
frame_pwm_obj_group_bin_0303 = frame (4k)
frame_pwm_obj_group_bin_0304 = frame (4k)
frame_pwm_obj_group_bin_0305 = frame (4k)
frame_pwm_obj_group_bin_0306 = frame (4k)
frame_pwm_obj_group_bin_0307 = frame (4k)
frame_pwm_obj_group_bin_0308 = frame (4k)
frame_pwm_obj_group_bin_0309 = frame (4k)
frame_pwm_obj_group_bin_0310 = frame (4k)
frame_pwm_obj_group_bin_0311 = frame (4k)
frame_pwm_obj_group_bin_0312 = frame (4k)
frame_pwm_obj_group_bin_0314 = frame (4k)
frame_pwm_obj_group_bin_0315 = frame (4k)
frame_pwm_obj_group_bin_0316 = frame (4k)
frame_pwm_obj_group_bin_0317 = frame (4k)
frame_pwm_obj_group_bin_0318 = frame (4k)
frame_pwm_obj_group_bin_0319 = frame (4k)
frame_pwm_obj_group_bin_0320 = frame (4k)
frame_pwm_obj_group_bin_0321 = frame (4k)
frame_pwm_obj_group_bin_0322 = frame (4k)
frame_pwm_obj_group_bin_0323 = frame (4k)
frame_pwm_obj_group_bin_0324 = frame (4k)
frame_pwm_obj_group_bin_0325 = frame (4k)
frame_pwm_obj_group_bin_0326 = frame (4k)
frame_pwm_obj_group_bin_0327 = frame (4k)
frame_pwm_obj_group_bin_0328 = frame (4k)
frame_pwm_obj_group_bin_0329 = frame (4k)
frame_pwm_obj_group_bin_0330 = frame (4k)
frame_pwm_obj_group_bin_0331 = frame (4k)
frame_pwm_obj_group_bin_0332 = frame (4k)
frame_pwm_obj_group_bin_0333 = frame (4k)
frame_pwm_obj_group_bin_0334 = frame (4k)
frame_spi_obj_group_bin_0000 = frame (4k)
frame_spi_obj_group_bin_0001 = frame (4k)
frame_spi_obj_group_bin_0002 = frame (4k)
frame_spi_obj_group_bin_0003 = frame (4k)
frame_spi_obj_group_bin_0004 = frame (4k)
frame_spi_obj_group_bin_0005 = frame (4k)
frame_spi_obj_group_bin_0006 = frame (4k)
frame_spi_obj_group_bin_0007 = frame (4k)
frame_spi_obj_group_bin_0008 = frame (4k)
frame_spi_obj_group_bin_0010 = frame (4k)
frame_spi_obj_group_bin_0011 = frame (4k)
frame_spi_obj_group_bin_0012 = frame (4k)
frame_spi_obj_group_bin_0013 = frame (4k)
frame_spi_obj_group_bin_0014 = frame (4k)
frame_spi_obj_group_bin_0015 = frame (4k)
frame_spi_obj_group_bin_0016 = frame (4k)
frame_spi_obj_group_bin_0017 = frame (4k)
frame_spi_obj_group_bin_0018 = frame (4k)
frame_spi_obj_group_bin_0019 = frame (4k)
frame_spi_obj_group_bin_0020 = frame (4k)
frame_spi_obj_group_bin_0021 = frame (4k)
frame_spi_obj_group_bin_0022 = frame (4k)
frame_spi_obj_group_bin_0023 = frame (4k)
frame_spi_obj_group_bin_0024 = frame (4k)
frame_spi_obj_group_bin_0025 = frame (4k)
frame_spi_obj_group_bin_0026 = frame (4k)
frame_spi_obj_group_bin_0027 = frame (4k)
frame_spi_obj_group_bin_0028 = frame (4k)
frame_spi_obj_group_bin_0029 = frame (4k)
frame_spi_obj_group_bin_0030 = frame (4k)
frame_spi_obj_group_bin_0031 = frame (4k)
frame_spi_obj_group_bin_0032 = frame (4k)
frame_spi_obj_group_bin_0033 = frame (4k)
frame_spi_obj_group_bin_0034 = frame (4k)
frame_spi_obj_group_bin_0035 = frame (4k)
frame_spi_obj_group_bin_0036 = frame (4k)
frame_spi_obj_group_bin_0037 = frame (4k)
frame_spi_obj_group_bin_0038 = frame (4k)
frame_spi_obj_group_bin_0039 = frame (4k)
frame_spi_obj_group_bin_0040 = frame (4k)
frame_spi_obj_group_bin_0041 = frame (4k)
frame_spi_obj_group_bin_0042 = frame (4k)
frame_spi_obj_group_bin_0043 = frame (4k)
frame_spi_obj_group_bin_0044 = frame (4k)
frame_spi_obj_group_bin_0045 = frame (4k)
frame_spi_obj_group_bin_0046 = frame (4k)
frame_spi_obj_group_bin_0047 = frame (4k)
frame_spi_obj_group_bin_0048 = frame (4k)
frame_spi_obj_group_bin_0049 = frame (4k)
frame_spi_obj_group_bin_0050 = frame (4k)
frame_spi_obj_group_bin_0051 = frame (4k)
frame_spi_obj_group_bin_0052 = frame (4k)
frame_spi_obj_group_bin_0053 = frame (4k)
frame_spi_obj_group_bin_0054 = frame (4k)
frame_spi_obj_group_bin_0055 = frame (4k)
frame_spi_obj_group_bin_0056 = frame (4k)
frame_spi_obj_group_bin_0057 = frame (4k)
frame_spi_obj_group_bin_0059 = frame (4k)
frame_spi_obj_group_bin_0060 = frame (4k)
frame_spi_obj_group_bin_0061 = frame (4k)
frame_spi_obj_group_bin_0062 = frame (4k)
frame_spi_obj_group_bin_0064 = frame (4k)
frame_spi_obj_group_bin_0065 = frame (4k)
frame_spi_obj_group_bin_0066 = frame (4k)
frame_spi_obj_group_bin_0067 = frame (4k)
frame_spi_obj_group_bin_0068 = frame (4k)
frame_spi_obj_group_bin_0069 = frame (4k)
frame_spi_obj_group_bin_0070 = frame (4k)
frame_spi_obj_group_bin_0071 = frame (4k)
frame_spi_obj_group_bin_0072 = frame (4k)
frame_spi_obj_group_bin_0073 = frame (4k)
frame_spi_obj_group_bin_0074 = frame (4k)
frame_spi_obj_group_bin_0075 = frame (4k)
frame_spi_obj_group_bin_0076 = frame (4k)
frame_spi_obj_group_bin_0077 = frame (4k)
frame_spi_obj_group_bin_0078 = frame (4k)
frame_spi_obj_group_bin_0079 = frame (4k)
frame_spi_obj_group_bin_0080 = frame (4k)
frame_spi_obj_group_bin_0081 = frame (4k)
frame_spi_obj_group_bin_0082 = frame (4k)
frame_spi_obj_group_bin_0083 = frame (4k)
frame_spi_obj_group_bin_0084 = frame (4k)
frame_spi_obj_group_bin_0085 = frame (4k)
frame_spi_obj_group_bin_0086 = frame (4k)
frame_spi_obj_group_bin_0087 = frame (4k)
frame_spi_obj_group_bin_0088 = frame (4k)
frame_spi_obj_group_bin_0089 = frame (4k)
frame_spi_obj_group_bin_0090 = frame (4k)
frame_spi_obj_group_bin_0091 = frame (4k)
frame_spi_obj_group_bin_0092 = frame (4k)
frame_spi_obj_group_bin_0093 = frame (4k)
frame_spi_obj_group_bin_0094 = frame (4k)
frame_spi_obj_group_bin_0095 = frame (4k)
frame_spi_obj_group_bin_0097 = frame (4k)
frame_spi_obj_group_bin_0098 = frame (4k)
frame_spi_obj_group_bin_0099 = frame (4k)
frame_spi_obj_group_bin_0100 = frame (4k)
frame_spi_obj_group_bin_0101 = frame (4k)
frame_spi_obj_group_bin_0102 = frame (4k)
frame_spi_obj_group_bin_0103 = frame (4k)
frame_spi_obj_group_bin_0104 = frame (4k)
frame_spi_obj_group_bin_0105 = frame (4k)
frame_spi_obj_group_bin_0106 = frame (4k)
frame_spi_obj_group_bin_0107 = frame (4k)
frame_spi_obj_group_bin_0109 = frame (4k)
frame_spi_obj_group_bin_0110 = frame (4k)
frame_spi_obj_group_bin_0111 = frame (4k)
frame_spi_obj_group_bin_0112 = frame (4k)
frame_spi_obj_group_bin_0113 = frame (4k)
frame_spi_obj_group_bin_0114 = frame (4k)
frame_spi_obj_group_bin_0115 = frame (4k)
frame_spi_obj_group_bin_0116 = frame (4k)
frame_spi_obj_group_bin_0117 = frame (4k)
frame_spi_obj_group_bin_0118 = frame (4k)
frame_spi_obj_group_bin_0119 = frame (4k)
frame_spi_obj_group_bin_0120 = frame (4k)
frame_spi_obj_group_bin_0121 = frame (4k)
frame_spi_obj_group_bin_0122 = frame (4k)
frame_spi_obj_group_bin_0123 = frame (4k)
frame_spi_obj_group_bin_0124 = frame (4k)
frame_spi_obj_group_bin_0125 = frame (4k)
frame_spi_obj_group_bin_0126 = frame (4k)
frame_spi_obj_group_bin_0127 = frame (4k)
frame_spi_obj_group_bin_0128 = frame (4k)
frame_spi_obj_group_bin_0129 = frame (4k)
frame_spi_obj_group_bin_0130 = frame (4k)
frame_spi_obj_group_bin_0131 = frame (4k)
frame_spi_obj_group_bin_0132 = frame (4k)
frame_spi_obj_group_bin_0133 = frame (4k)
frame_spi_obj_group_bin_0134 = frame (4k)
frame_spi_obj_group_bin_0135 = frame (4k)
frame_spi_obj_group_bin_0136 = frame (4k)
frame_spi_obj_group_bin_0137 = frame (4k)
frame_spi_obj_group_bin_0138 = frame (4k)
frame_spi_obj_group_bin_0139 = frame (4k)
frame_spi_obj_group_bin_0140 = frame (4k)
frame_spi_obj_group_bin_0141 = frame (4k)
frame_spi_obj_group_bin_0142 = frame (4k)
frame_spi_obj_group_bin_0143 = frame (4k)
frame_spi_obj_group_bin_0145 = frame (4k)
frame_spi_obj_group_bin_0146 = frame (4k)
frame_spi_obj_group_bin_0147 = frame (4k)
frame_spi_obj_group_bin_0148 = frame (4k)
frame_spi_obj_group_bin_0149 = frame (4k)
frame_spi_obj_group_bin_0150 = frame (4k)
frame_spi_obj_group_bin_0151 = frame (4k)
frame_spi_obj_group_bin_0152 = frame (4k)
frame_spi_obj_group_bin_0153 = frame (4k)
frame_spi_obj_group_bin_0154 = frame (4k)
frame_spi_obj_group_bin_0155 = frame (4k)
frame_spi_obj_group_bin_0156 = frame (4k)
frame_spi_obj_group_bin_0157 = frame (4k)
frame_spi_obj_group_bin_0158 = frame (4k)
frame_spi_obj_group_bin_0159 = frame (4k)
frame_spi_obj_group_bin_0160 = frame (4k)
frame_spi_obj_group_bin_0161 = frame (4k)
frame_spi_obj_group_bin_0162 = frame (4k)
frame_spi_obj_group_bin_0163 = frame (4k)
frame_spi_obj_group_bin_0164 = frame (4k)
frame_spi_obj_group_bin_0165 = frame (4k)
frame_spi_obj_group_bin_0166 = frame (4k)
frame_spi_obj_group_bin_0167 = frame (4k)
frame_spi_obj_group_bin_0168 = frame (4k)
frame_spi_obj_group_bin_0169 = frame (4k)
frame_spi_obj_group_bin_0170 = frame (4k)
frame_spi_obj_group_bin_0171 = frame (4k)
frame_spi_obj_group_bin_0172 = frame (4k)
frame_spi_obj_group_bin_0173 = frame (4k)
frame_spi_obj_group_bin_0174 = frame (4k)
frame_spi_obj_group_bin_0175 = frame (4k)
frame_spi_obj_group_bin_0176 = frame (4k)
frame_spi_obj_group_bin_0177 = frame (4k)
frame_spi_obj_group_bin_0178 = frame (4k)
frame_spi_obj_group_bin_0179 = frame (4k)
frame_spi_obj_group_bin_0180 = frame (4k)
frame_spi_obj_group_bin_0181 = frame (4k)
frame_spi_obj_group_bin_0182 = frame (4k)
frame_spi_obj_group_bin_0183 = frame (4k)
frame_spi_obj_group_bin_0184 = frame (4k)
frame_spi_obj_group_bin_0185 = frame (4k)
frame_spi_obj_group_bin_0186 = frame (4k)
frame_spi_obj_group_bin_0187 = frame (4k)
frame_spi_obj_group_bin_0189 = frame (4k)
frame_spi_obj_group_bin_0190 = frame (4k)
frame_spi_obj_group_bin_0191 = frame (4k)
frame_spi_obj_group_bin_0192 = frame (4k)
frame_spi_obj_group_bin_0193 = frame (4k)
frame_spi_obj_group_bin_0194 = frame (4k)
frame_spi_obj_group_bin_0195 = frame (4k)
frame_spi_obj_group_bin_0196 = frame (4k)
frame_spi_obj_group_bin_0197 = frame (4k)
frame_spi_obj_group_bin_0198 = frame (4k)
frame_spi_obj_group_bin_0199 = frame (4k)
frame_spi_obj_group_bin_0200 = frame (4k)
frame_spi_obj_group_bin_0201 = frame (4k)
frame_spi_obj_group_bin_0203 = frame (4k)
frame_spi_obj_group_bin_0204 = frame (4k)
frame_spi_obj_group_bin_0205 = frame (4k)
frame_spi_obj_group_bin_0207 = frame (4k)
frame_spi_obj_group_bin_0208 = frame (4k)
frame_spi_obj_group_bin_0209 = frame (4k)
frame_spi_obj_group_bin_0210 = frame (4k)
frame_spi_obj_group_bin_0211 = frame (4k)
frame_spi_obj_group_bin_0212 = frame (4k)
frame_spi_obj_group_bin_0213 = frame (4k)
frame_spi_obj_group_bin_0214 = frame (4k)
frame_spi_obj_group_bin_0215 = frame (4k)
frame_spi_obj_group_bin_0216 = frame (4k)
frame_spi_obj_group_bin_0217 = frame (4k)
frame_spi_obj_group_bin_0218 = frame (4k)
frame_spi_obj_group_bin_0219 = frame (4k)
frame_spi_obj_group_bin_0220 = frame (4k)
frame_spi_obj_group_bin_0221 = frame (4k)
frame_spi_obj_group_bin_0222 = frame (4k)
frame_spi_obj_group_bin_0223 = frame (4k)
frame_spi_obj_group_bin_0224 = frame (4k)
frame_spi_obj_group_bin_0225 = frame (4k)
frame_spi_obj_group_bin_0226 = frame (4k)
frame_spi_obj_group_bin_0227 = frame (4k)
frame_spi_obj_group_bin_0228 = frame (4k)
frame_spi_obj_group_bin_0229 = frame (4k)
frame_spi_obj_group_bin_0231 = frame (4k)
frame_spi_obj_group_bin_0232 = frame (4k)
frame_spi_obj_group_bin_0233 = frame (4k)
frame_spi_obj_group_bin_0234 = frame (4k)
frame_spi_obj_group_bin_0235 = frame (4k)
frame_spi_obj_group_bin_0236 = frame (4k)
frame_spi_obj_group_bin_0237 = frame (4k)
frame_spi_obj_group_bin_0238 = frame (4k)
frame_spi_obj_group_bin_0239 = frame (4k)
frame_spi_obj_group_bin_0240 = frame (4k)
frame_spi_obj_group_bin_0241 = frame (4k)
frame_spi_obj_group_bin_0242 = frame (4k)
frame_spi_obj_group_bin_0243 = frame (4k)
frame_spi_obj_group_bin_0244 = frame (4k)
frame_spi_obj_group_bin_0245 = frame (4k)
frame_spi_obj_group_bin_0246 = frame (4k, paddr: 0x12d30000)
frame_spi_obj_group_bin_0247 = frame (4k)
frame_spi_obj_group_bin_0248 = frame (4k)
frame_spi_obj_group_bin_0249 = frame (4k)
frame_spi_obj_group_bin_0250 = frame (4k)
frame_spi_obj_group_bin_0251 = frame (4k)
frame_spi_obj_group_bin_0252 = frame (4k)
frame_spi_obj_group_bin_0253 = frame (4k)
frame_spi_obj_group_bin_0254 = frame (4k)
frame_spi_obj_group_bin_0255 = frame (4k)
frame_spi_obj_group_bin_0256 = frame (4k)
frame_spi_obj_group_bin_0257 = frame (4k)
frame_spi_obj_group_bin_0258 = frame (4k)
frame_spi_obj_group_bin_0259 = frame (4k)
frame_spi_obj_group_bin_0261 = frame (4k)
frame_spi_obj_group_bin_0262 = frame (4k)
frame_spi_obj_group_bin_0263 = frame (4k)
frame_spi_obj_group_bin_0264 = frame (4k)
frame_spi_obj_group_bin_0265 = frame (4k)
frame_spi_obj_group_bin_0266 = frame (4k)
frame_spi_obj_group_bin_0267 = frame (4k)
frame_spi_obj_group_bin_0268 = frame (4k)
frame_spi_obj_group_bin_0270 = frame (4k)
frame_spi_obj_group_bin_0271 = frame (4k)
frame_spi_obj_group_bin_0273 = frame (4k)
frame_spi_obj_group_bin_0274 = frame (4k)
frame_spi_obj_group_bin_0275 = frame (4k)
frame_spi_obj_group_bin_0276 = frame (4k)
frame_spi_obj_group_bin_0277 = frame (4k)
frame_spi_obj_group_bin_0278 = frame (4k)
frame_spi_obj_group_bin_0279 = frame (4k)
frame_spi_obj_group_bin_0280 = frame (4k)
frame_spi_obj_group_bin_0281 = frame (4k)
frame_spi_obj_group_bin_0282 = frame (4k)
frame_spi_obj_group_bin_0283 = frame (4k)
frame_spi_obj_group_bin_0284 = frame (4k)
frame_spi_obj_group_bin_0285 = frame (4k)
frame_spi_obj_group_bin_0286 = frame (4k)
frame_spi_obj_group_bin_0288 = frame (4k)
frame_spi_obj_group_bin_0290 = frame (4k)
frame_spi_obj_group_bin_0292 = frame (4k)
frame_spi_obj_group_bin_0293 = frame (4k)
frame_spi_obj_group_bin_0294 = frame (4k)
frame_spi_obj_group_bin_0295 = frame (4k)
frame_spi_obj_group_bin_0296 = frame (4k)
frame_spi_obj_group_bin_0298 = frame (4k)
frame_spi_obj_group_bin_0299 = frame (4k)
frame_spi_obj_group_bin_0300 = frame (4k)
frame_spi_obj_group_bin_0301 = frame (4k)
frame_spi_obj_group_bin_0302 = frame (4k)
frame_spi_obj_group_bin_0303 = frame (4k)
frame_spi_obj_group_bin_0304 = frame (4k)
frame_spi_obj_group_bin_0305 = frame (4k)
frame_spi_obj_group_bin_0306 = frame (4k)
frame_spi_obj_group_bin_0307 = frame (4k)
frame_spi_obj_group_bin_0308 = frame (4k)
frame_spi_obj_group_bin_0309 = frame (4k)
frame_spi_obj_group_bin_0310 = frame (4k)
frame_spi_obj_group_bin_0311 = frame (4k)
frame_spi_obj_group_bin_0312 = frame (4k)
frame_spi_obj_group_bin_0313 = frame (4k)
frame_spi_obj_group_bin_0314 = frame (4k)
frame_spi_obj_group_bin_0315 = frame (4k)
frame_spi_obj_group_bin_0316 = frame (4k)
frame_timer_obj_group_bin_0000 = frame (4k)
frame_timer_obj_group_bin_0001 = frame (4k)
frame_timer_obj_group_bin_0002 = frame (4k)
frame_timer_obj_group_bin_0003 = frame (4k)
frame_timer_obj_group_bin_0004 = frame (4k)
frame_timer_obj_group_bin_0005 = frame (4k)
frame_timer_obj_group_bin_0006 = frame (4k)
frame_timer_obj_group_bin_0007 = frame (4k)
frame_timer_obj_group_bin_0008 = frame (4k)
frame_timer_obj_group_bin_0009 = frame (4k)
frame_timer_obj_group_bin_0010 = frame (4k)
frame_timer_obj_group_bin_0011 = frame (4k)
frame_timer_obj_group_bin_0012 = frame (4k)
frame_timer_obj_group_bin_0013 = frame (4k)
frame_timer_obj_group_bin_0014 = frame (4k)
frame_timer_obj_group_bin_0016 = frame (4k)
frame_timer_obj_group_bin_0017 = frame (4k)
frame_timer_obj_group_bin_0018 = frame (4k)
frame_timer_obj_group_bin_0019 = frame (4k)
frame_timer_obj_group_bin_0020 = frame (4k)
frame_timer_obj_group_bin_0021 = frame (4k)
frame_timer_obj_group_bin_0022 = frame (4k)
frame_timer_obj_group_bin_0023 = frame (4k)
frame_timer_obj_group_bin_0024 = frame (4k)
frame_timer_obj_group_bin_0025 = frame (4k)
frame_timer_obj_group_bin_0026 = frame (4k)
frame_timer_obj_group_bin_0027 = frame (4k)
frame_timer_obj_group_bin_0028 = frame (4k)
frame_timer_obj_group_bin_0029 = frame (4k)
frame_timer_obj_group_bin_0030 = frame (4k)
frame_timer_obj_group_bin_0031 = frame (4k)
frame_timer_obj_group_bin_0032 = frame (4k)
frame_timer_obj_group_bin_0033 = frame (4k)
frame_timer_obj_group_bin_0034 = frame (4k)
frame_timer_obj_group_bin_0035 = frame (4k)
frame_timer_obj_group_bin_0036 = frame (4k)
frame_timer_obj_group_bin_0037 = frame (4k)
frame_timer_obj_group_bin_0038 = frame (4k)
frame_timer_obj_group_bin_0039 = frame (4k)
frame_timer_obj_group_bin_0040 = frame (4k)
frame_timer_obj_group_bin_0041 = frame (4k)
frame_timer_obj_group_bin_0042 = frame (4k)
frame_timer_obj_group_bin_0043 = frame (4k)
frame_timer_obj_group_bin_0044 = frame (4k)
frame_timer_obj_group_bin_0045 = frame (4k)
frame_timer_obj_group_bin_0046 = frame (4k)
frame_timer_obj_group_bin_0047 = frame (4k)
frame_timer_obj_group_bin_0048 = frame (4k)
frame_timer_obj_group_bin_0049 = frame (4k)
frame_timer_obj_group_bin_0050 = frame (4k)
frame_timer_obj_group_bin_0051 = frame (4k)
frame_timer_obj_group_bin_0052 = frame (4k)
frame_timer_obj_group_bin_0053 = frame (4k)
frame_timer_obj_group_bin_0054 = frame (4k)
frame_timer_obj_group_bin_0055 = frame (4k)
frame_timer_obj_group_bin_0056 = frame (4k)
frame_timer_obj_group_bin_0057 = frame (4k)
frame_timer_obj_group_bin_0058 = frame (4k)
frame_timer_obj_group_bin_0059 = frame (4k)
frame_timer_obj_group_bin_0060 = frame (4k)
frame_timer_obj_group_bin_0061 = frame (4k)
frame_timer_obj_group_bin_0062 = frame (4k)
frame_timer_obj_group_bin_0063 = frame (4k)
frame_timer_obj_group_bin_0064 = frame (4k)
frame_timer_obj_group_bin_0065 = frame (4k)
frame_timer_obj_group_bin_0066 = frame (4k)
frame_timer_obj_group_bin_0067 = frame (4k)
frame_timer_obj_group_bin_0068 = frame (4k)
frame_timer_obj_group_bin_0069 = frame (4k)
frame_timer_obj_group_bin_0070 = frame (4k)
frame_timer_obj_group_bin_0071 = frame (4k)
frame_timer_obj_group_bin_0072 = frame (4k)
frame_timer_obj_group_bin_0073 = frame (4k)
frame_timer_obj_group_bin_0074 = frame (4k)
frame_timer_obj_group_bin_0075 = frame (4k)
frame_timer_obj_group_bin_0077 = frame (4k)
frame_timer_obj_group_bin_0078 = frame (4k)
frame_timer_obj_group_bin_0079 = frame (4k)
frame_timer_obj_group_bin_0080 = frame (4k)
frame_timer_obj_group_bin_0081 = frame (4k)
frame_timer_obj_group_bin_0082 = frame (4k)
frame_timer_obj_group_bin_0083 = frame (4k)
frame_timer_obj_group_bin_0084 = frame (4k)
frame_timer_obj_group_bin_0085 = frame (4k)
frame_timer_obj_group_bin_0086 = frame (4k)
frame_timer_obj_group_bin_0087 = frame (4k)
frame_timer_obj_group_bin_0088 = frame (4k)
frame_timer_obj_group_bin_0089 = frame (4k)
frame_timer_obj_group_bin_0090 = frame (4k)
frame_timer_obj_group_bin_0091 = frame (4k)
frame_timer_obj_group_bin_0092 = frame (4k)
frame_timer_obj_group_bin_0093 = frame (4k)
frame_timer_obj_group_bin_0094 = frame (4k)
frame_timer_obj_group_bin_0095 = frame (4k)
frame_timer_obj_group_bin_0096 = frame (4k)
frame_timer_obj_group_bin_0097 = frame (4k)
frame_timer_obj_group_bin_0098 = frame (4k)
frame_timer_obj_group_bin_0100 = frame (4k)
frame_timer_obj_group_bin_0101 = frame (4k)
frame_timer_obj_group_bin_0102 = frame (4k)
frame_timer_obj_group_bin_0103 = frame (4k)
frame_timer_obj_group_bin_0104 = frame (4k)
frame_timer_obj_group_bin_0105 = frame (4k)
frame_timer_obj_group_bin_0106 = frame (4k)
frame_timer_obj_group_bin_0107 = frame (4k)
frame_timer_obj_group_bin_0108 = frame (4k)
frame_timer_obj_group_bin_0109 = frame (4k)
frame_timer_obj_group_bin_0110 = frame (4k)
frame_timer_obj_group_bin_0111 = frame (4k)
frame_timer_obj_group_bin_0112 = frame (4k)
frame_timer_obj_group_bin_0113 = frame (4k)
frame_timer_obj_group_bin_0114 = frame (4k)
frame_timer_obj_group_bin_0115 = frame (4k)
frame_timer_obj_group_bin_0116 = frame (4k)
frame_timer_obj_group_bin_0117 = frame (4k)
frame_timer_obj_group_bin_0118 = frame (4k)
frame_timer_obj_group_bin_0119 = frame (4k)
frame_timer_obj_group_bin_0120 = frame (4k)
frame_timer_obj_group_bin_0122 = frame (4k)
frame_timer_obj_group_bin_0123 = frame (4k)
frame_timer_obj_group_bin_0124 = frame (4k)
frame_timer_obj_group_bin_0125 = frame (4k)
frame_timer_obj_group_bin_0126 = frame (4k)
frame_timer_obj_group_bin_0127 = frame (4k)
frame_timer_obj_group_bin_0128 = frame (4k)
frame_timer_obj_group_bin_0129 = frame (4k)
frame_timer_obj_group_bin_0130 = frame (4k)
frame_timer_obj_group_bin_0131 = frame (4k)
frame_timer_obj_group_bin_0132 = frame (4k)
frame_timer_obj_group_bin_0133 = frame (4k)
frame_timer_obj_group_bin_0134 = frame (4k)
frame_timer_obj_group_bin_0135 = frame (4k)
frame_timer_obj_group_bin_0136 = frame (4k)
frame_timer_obj_group_bin_0138 = frame (4k)
frame_timer_obj_group_bin_0139 = frame (4k)
frame_timer_obj_group_bin_0140 = frame (4k)
frame_timer_obj_group_bin_0141 = frame (4k)
frame_timer_obj_group_bin_0142 = frame (4k)
frame_timer_obj_group_bin_0143 = frame (4k)
frame_timer_obj_group_bin_0144 = frame (4k)
frame_timer_obj_group_bin_0145 = frame (4k)
frame_timer_obj_group_bin_0146 = frame (4k)
frame_timer_obj_group_bin_0147 = frame (4k)
frame_timer_obj_group_bin_0148 = frame (4k)
frame_timer_obj_group_bin_0149 = frame (4k)
frame_timer_obj_group_bin_0150 = frame (4k)
frame_timer_obj_group_bin_0151 = frame (4k)
frame_timer_obj_group_bin_0153 = frame (4k)
frame_timer_obj_group_bin_0154 = frame (4k)
frame_timer_obj_group_bin_0155 = frame (4k)
frame_timer_obj_group_bin_0156 = frame (4k)
frame_timer_obj_group_bin_0157 = frame (4k)
frame_timer_obj_group_bin_0158 = frame (4k)
frame_timer_obj_group_bin_0159 = frame (4k)
frame_timer_obj_group_bin_0160 = frame (4k)
frame_timer_obj_group_bin_0161 = frame (4k)
frame_timer_obj_group_bin_0162 = frame (4k)
frame_timer_obj_group_bin_0163 = frame (4k)
frame_timer_obj_group_bin_0164 = frame (4k)
frame_timer_obj_group_bin_0165 = frame (4k)
frame_timer_obj_group_bin_0166 = frame (4k)
frame_timer_obj_group_bin_0167 = frame (4k)
frame_timer_obj_group_bin_0168 = frame (4k)
frame_timer_obj_group_bin_0169 = frame (4k)
frame_timer_obj_group_bin_0170 = frame (4k)
frame_timer_obj_group_bin_0171 = frame (4k)
frame_timer_obj_group_bin_0172 = frame (4k)
frame_timer_obj_group_bin_0173 = frame (4k)
frame_timer_obj_group_bin_0174 = frame (4k)
frame_timer_obj_group_bin_0175 = frame (4k)
frame_timer_obj_group_bin_0176 = frame (4k)
frame_timer_obj_group_bin_0178 = frame (4k)
frame_timer_obj_group_bin_0179 = frame (4k)
frame_timer_obj_group_bin_0180 = frame (4k)
frame_timer_obj_group_bin_0181 = frame (4k)
frame_timer_obj_group_bin_0182 = frame (4k)
frame_timer_obj_group_bin_0183 = frame (4k)
frame_timer_obj_group_bin_0185 = frame (4k)
frame_timer_obj_group_bin_0186 = frame (4k)
frame_timer_obj_group_bin_0187 = frame (4k)
frame_timer_obj_group_bin_0188 = frame (4k)
frame_timer_obj_group_bin_0189 = frame (4k)
frame_timer_obj_group_bin_0190 = frame (4k)
frame_timer_obj_group_bin_0191 = frame (4k)
frame_timer_obj_group_bin_0192 = frame (4k)
frame_timer_obj_group_bin_0193 = frame (4k)
frame_timer_obj_group_bin_0194 = frame (4k)
frame_timer_obj_group_bin_0195 = frame (4k)
frame_timer_obj_group_bin_0196 = frame (4k)
frame_timer_obj_group_bin_0197 = frame (4k)
frame_timer_obj_group_bin_0198 = frame (4k)
frame_timer_obj_group_bin_0199 = frame (4k)
frame_timer_obj_group_bin_0200 = frame (4k)
frame_timer_obj_group_bin_0201 = frame (4k)
frame_timer_obj_group_bin_0202 = frame (4k)
frame_timer_obj_group_bin_0203 = frame (4k)
frame_timer_obj_group_bin_0204 = frame (4k)
frame_timer_obj_group_bin_0205 = frame (4k)
frame_timer_obj_group_bin_0206 = frame (4k)
frame_timer_obj_group_bin_0207 = frame (4k)
frame_timer_obj_group_bin_0208 = frame (4k)
frame_timer_obj_group_bin_0209 = frame (4k)
frame_timer_obj_group_bin_0210 = frame (4k)
frame_timer_obj_group_bin_0211 = frame (4k)
frame_timer_obj_group_bin_0212 = frame (4k)
frame_timer_obj_group_bin_0213 = frame (4k)
frame_timer_obj_group_bin_0214 = frame (4k)
frame_timer_obj_group_bin_0215 = frame (4k)
frame_timer_obj_group_bin_0216 = frame (4k)
frame_timer_obj_group_bin_0217 = frame (4k)
frame_timer_obj_group_bin_0219 = frame (4k)
frame_timer_obj_group_bin_0220 = frame (4k)
frame_timer_obj_group_bin_0221 = frame (4k)
frame_timer_obj_group_bin_0222 = frame (4k)
frame_timer_obj_group_bin_0223 = frame (4k)
frame_timer_obj_group_bin_0224 = frame (4k)
frame_timer_obj_group_bin_0225 = frame (4k)
frame_timer_obj_group_bin_0226 = frame (4k)
frame_timer_obj_group_bin_0227 = frame (4k)
frame_timer_obj_group_bin_0228 = frame (4k)
frame_timer_obj_group_bin_0229 = frame (4k)
frame_timer_obj_group_bin_0230 = frame (4k)
frame_timer_obj_group_bin_0231 = frame (4k)
frame_timer_obj_group_bin_0232 = frame (4k)
frame_timer_obj_group_bin_0233 = frame (4k)
frame_timer_obj_group_bin_0234 = frame (4k, paddr: 0x12dd0000)
frame_timer_obj_group_bin_0235 = frame (4k)
frame_timer_obj_group_bin_0236 = frame (4k)
frame_timer_obj_group_bin_0237 = frame (4k)
frame_timer_obj_group_bin_0238 = frame (4k)
frame_timer_obj_group_bin_0239 = frame (4k)
frame_timer_obj_group_bin_0240 = frame (4k)
frame_timer_obj_group_bin_0241 = frame (4k)
frame_timer_obj_group_bin_0242 = frame (4k)
frame_timer_obj_group_bin_0243 = frame (4k)
frame_timer_obj_group_bin_0244 = frame (4k)
frame_timer_obj_group_bin_0245 = frame (4k)
frame_timer_obj_group_bin_0246 = frame (4k)
frame_timer_obj_group_bin_0248 = frame (4k)
frame_timer_obj_group_bin_0250 = frame (4k)
frame_timer_obj_group_bin_0251 = frame (4k)
frame_timer_obj_group_bin_0252 = frame (4k)
frame_timer_obj_group_bin_0253 = frame (4k)
frame_timer_obj_group_bin_0254 = frame (4k)
frame_timer_obj_group_bin_0255 = frame (4k)
frame_timer_obj_group_bin_0257 = frame (4k)
frame_timer_obj_group_bin_0258 = frame (4k)
frame_timer_obj_group_bin_0259 = frame (4k)
frame_timer_obj_group_bin_0260 = frame (4k)
frame_timer_obj_group_bin_0261 = frame (4k)
frame_timer_obj_group_bin_0262 = frame (4k)
frame_timer_obj_group_bin_0263 = frame (4k)
frame_timer_obj_group_bin_0264 = frame (4k)
frame_timer_obj_group_bin_0265 = frame (4k)
frame_timer_obj_group_bin_0266 = frame (4k)
frame_timer_obj_group_bin_0267 = frame (4k)
frame_timer_obj_group_bin_0268 = frame (4k)
frame_timer_obj_group_bin_0269 = frame (4k)
frame_timer_obj_group_bin_0270 = frame (4k)
frame_timer_obj_group_bin_0271 = frame (4k)
frame_timer_obj_group_bin_0272 = frame (4k)
frame_timer_obj_group_bin_0273 = frame (4k)
frame_timer_obj_group_bin_0274 = frame (4k)
frame_timer_obj_group_bin_0275 = frame (4k)
frame_timer_obj_group_bin_0276 = frame (4k)
frame_timer_obj_group_bin_0277 = frame (4k)
frame_timer_obj_group_bin_0278 = frame (4k)
frame_timer_obj_group_bin_0279 = frame (4k)
frame_timer_obj_group_bin_0280 = frame (4k)
frame_timer_obj_group_bin_0281 = frame (4k)
frame_timer_obj_group_bin_0282 = frame (4k)
frame_timer_obj_group_bin_0283 = frame (4k)
frame_timer_obj_group_bin_0284 = frame (4k)
frame_timer_obj_group_bin_0285 = frame (4k)
frame_timer_obj_group_bin_0286 = frame (4k)
frame_timer_obj_group_bin_0287 = frame (4k)
frame_timer_obj_group_bin_0288 = frame (4k)
frame_timer_obj_group_bin_0289 = frame (4k)
frame_timer_obj_group_bin_0290 = frame (4k)
frame_timer_obj_group_bin_0291 = frame (4k)
frame_timer_obj_group_bin_0292 = frame (4k)
frame_timer_obj_group_bin_0293 = frame (4k)
frame_timer_obj_group_bin_0294 = frame (4k)
frame_timer_obj_group_bin_0295 = frame (4k)
frame_timer_obj_group_bin_0296 = frame (4k)
frame_timer_obj_group_bin_0297 = frame (4k)
frame_timer_obj_group_bin_0298 = frame (4k)
frame_timer_obj_group_bin_0299 = frame (4k)
frame_timer_obj_group_bin_0300 = frame (4k)
frame_uart_gcs_group_bin_0000 = frame (4k)
frame_uart_gcs_group_bin_0001 = frame (4k)
frame_uart_gcs_group_bin_0002 = frame (4k)
frame_uart_gcs_group_bin_0003 = frame (4k)
frame_uart_gcs_group_bin_0004 = frame (4k)
frame_uart_gcs_group_bin_0005 = frame (4k)
frame_uart_gcs_group_bin_0006 = frame (4k)
frame_uart_gcs_group_bin_0007 = frame (4k)
frame_uart_gcs_group_bin_0008 = frame (4k)
frame_uart_gcs_group_bin_0009 = frame (4k)
frame_uart_gcs_group_bin_0010 = frame (4k)
frame_uart_gcs_group_bin_0011 = frame (4k)
frame_uart_gcs_group_bin_0012 = frame (4k)
frame_uart_gcs_group_bin_0013 = frame (4k)
frame_uart_gcs_group_bin_0014 = frame (4k)
frame_uart_gcs_group_bin_0017 = frame (4k)
frame_uart_gcs_group_bin_0018 = frame (4k)
frame_uart_gcs_group_bin_0019 = frame (4k)
frame_uart_gcs_group_bin_0020 = frame (4k)
frame_uart_gcs_group_bin_0021 = frame (4k)
frame_uart_gcs_group_bin_0022 = frame (4k)
frame_uart_gcs_group_bin_0024 = frame (4k)
frame_uart_gcs_group_bin_0025 = frame (4k)
frame_uart_gcs_group_bin_0026 = frame (4k)
frame_uart_gcs_group_bin_0027 = frame (4k)
frame_uart_gcs_group_bin_0028 = frame (4k)
frame_uart_gcs_group_bin_0029 = frame (4k)
frame_uart_gcs_group_bin_0030 = frame (4k)
frame_uart_gcs_group_bin_0031 = frame (4k)
frame_uart_gcs_group_bin_0032 = frame (4k)
frame_uart_gcs_group_bin_0033 = frame (4k)
frame_uart_gcs_group_bin_0034 = frame (4k)
frame_uart_gcs_group_bin_0035 = frame (4k)
frame_uart_gcs_group_bin_0036 = frame (4k)
frame_uart_gcs_group_bin_0037 = frame (4k)
frame_uart_gcs_group_bin_0038 = frame (4k)
frame_uart_gcs_group_bin_0039 = frame (4k)
frame_uart_gcs_group_bin_0040 = frame (4k)
frame_uart_gcs_group_bin_0041 = frame (4k)
frame_uart_gcs_group_bin_0042 = frame (4k)
frame_uart_gcs_group_bin_0043 = frame (4k)
frame_uart_gcs_group_bin_0044 = frame (4k)
frame_uart_gcs_group_bin_0045 = frame (4k)
frame_uart_gcs_group_bin_0046 = frame (4k)
frame_uart_gcs_group_bin_0047 = frame (4k)
frame_uart_gcs_group_bin_0048 = frame (4k)
frame_uart_gcs_group_bin_0049 = frame (4k)
frame_uart_gcs_group_bin_0050 = frame (4k)
frame_uart_gcs_group_bin_0051 = frame (4k)
frame_uart_gcs_group_bin_0052 = frame (4k)
frame_uart_gcs_group_bin_0053 = frame (4k)
frame_uart_gcs_group_bin_0054 = frame (4k)
frame_uart_gcs_group_bin_0055 = frame (4k)
frame_uart_gcs_group_bin_0057 = frame (4k)
frame_uart_gcs_group_bin_0059 = frame (4k)
frame_uart_gcs_group_bin_0060 = frame (4k)
frame_uart_gcs_group_bin_0061 = frame (4k)
frame_uart_gcs_group_bin_0062 = frame (4k)
frame_uart_gcs_group_bin_0063 = frame (4k)
frame_uart_gcs_group_bin_0064 = frame (4k)
frame_uart_gcs_group_bin_0065 = frame (4k)
frame_uart_gcs_group_bin_0066 = frame (4k)
frame_uart_gcs_group_bin_0067 = frame (4k)
frame_uart_gcs_group_bin_0068 = frame (4k)
frame_uart_gcs_group_bin_0069 = frame (4k)
frame_uart_gcs_group_bin_0070 = frame (4k)
frame_uart_gcs_group_bin_0071 = frame (4k)
frame_uart_gcs_group_bin_0072 = frame (4k)
frame_uart_gcs_group_bin_0073 = frame (4k)
frame_uart_gcs_group_bin_0074 = frame (4k)
frame_uart_gcs_group_bin_0075 = frame (4k)
frame_uart_gcs_group_bin_0076 = frame (4k)
frame_uart_gcs_group_bin_0077 = frame (4k)
frame_uart_gcs_group_bin_0078 = frame (4k)
frame_uart_gcs_group_bin_0079 = frame (4k)
frame_uart_gcs_group_bin_0080 = frame (4k)
frame_uart_gcs_group_bin_0081 = frame (4k)
frame_uart_gcs_group_bin_0082 = frame (4k)
frame_uart_gcs_group_bin_0083 = frame (4k)
frame_uart_gcs_group_bin_0084 = frame (4k)
frame_uart_gcs_group_bin_0085 = frame (4k)
frame_uart_gcs_group_bin_0086 = frame (4k)
frame_uart_gcs_group_bin_0087 = frame (4k)
frame_uart_gcs_group_bin_0088 = frame (4k)
frame_uart_gcs_group_bin_0089 = frame (4k)
frame_uart_gcs_group_bin_0090 = frame (4k)
frame_uart_gcs_group_bin_0091 = frame (4k)
frame_uart_gcs_group_bin_0092 = frame (4k)
frame_uart_gcs_group_bin_0093 = frame (4k)
frame_uart_gcs_group_bin_0094 = frame (4k)
frame_uart_gcs_group_bin_0095 = frame (4k)
frame_uart_gcs_group_bin_0096 = frame (4k)
frame_uart_gcs_group_bin_0097 = frame (4k)
frame_uart_gcs_group_bin_0098 = frame (4k)
frame_uart_gcs_group_bin_0099 = frame (4k)
frame_uart_gcs_group_bin_0100 = frame (4k)
frame_uart_gcs_group_bin_0101 = frame (4k)
frame_uart_gcs_group_bin_0102 = frame (4k)
frame_uart_gcs_group_bin_0104 = frame (4k)
frame_uart_gcs_group_bin_0105 = frame (4k)
frame_uart_gcs_group_bin_0106 = frame (4k)
frame_uart_gcs_group_bin_0107 = frame (4k)
frame_uart_gcs_group_bin_0108 = frame (4k)
frame_uart_gcs_group_bin_0109 = frame (4k)
frame_uart_gcs_group_bin_0110 = frame (4k)
frame_uart_gcs_group_bin_0111 = frame (4k)
frame_uart_gcs_group_bin_0112 = frame (4k)
frame_uart_gcs_group_bin_0113 = frame (4k)
frame_uart_gcs_group_bin_0114 = frame (4k)
frame_uart_gcs_group_bin_0115 = frame (4k)
frame_uart_gcs_group_bin_0116 = frame (4k)
frame_uart_gcs_group_bin_0117 = frame (4k)
frame_uart_gcs_group_bin_0118 = frame (4k)
frame_uart_gcs_group_bin_0119 = frame (4k)
frame_uart_gcs_group_bin_0120 = frame (4k)
frame_uart_gcs_group_bin_0121 = frame (4k)
frame_uart_gcs_group_bin_0122 = frame (4k)
frame_uart_gcs_group_bin_0123 = frame (4k)
frame_uart_gcs_group_bin_0124 = frame (4k)
frame_uart_gcs_group_bin_0125 = frame (4k)
frame_uart_gcs_group_bin_0126 = frame (4k)
frame_uart_gcs_group_bin_0128 = frame (4k)
frame_uart_gcs_group_bin_0129 = frame (4k)
frame_uart_gcs_group_bin_0130 = frame (4k)
frame_uart_gcs_group_bin_0131 = frame (4k)
frame_uart_gcs_group_bin_0132 = frame (4k)
frame_uart_gcs_group_bin_0133 = frame (4k)
frame_uart_gcs_group_bin_0134 = frame (4k)
frame_uart_gcs_group_bin_0135 = frame (4k)
frame_uart_gcs_group_bin_0136 = frame (4k)
frame_uart_gcs_group_bin_0137 = frame (4k)
frame_uart_gcs_group_bin_0138 = frame (4k)
frame_uart_gcs_group_bin_0139 = frame (4k)
frame_uart_gcs_group_bin_0140 = frame (4k)
frame_uart_gcs_group_bin_0141 = frame (4k)
frame_uart_gcs_group_bin_0142 = frame (4k)
frame_uart_gcs_group_bin_0143 = frame (4k)
frame_uart_gcs_group_bin_0145 = frame (4k)
frame_uart_gcs_group_bin_0146 = frame (4k)
frame_uart_gcs_group_bin_0147 = frame (4k)
frame_uart_gcs_group_bin_0148 = frame (4k)
frame_uart_gcs_group_bin_0149 = frame (4k)
frame_uart_gcs_group_bin_0150 = frame (4k)
frame_uart_gcs_group_bin_0151 = frame (4k)
frame_uart_gcs_group_bin_0152 = frame (4k)
frame_uart_gcs_group_bin_0153 = frame (4k)
frame_uart_gcs_group_bin_0154 = frame (4k)
frame_uart_gcs_group_bin_0155 = frame (4k)
frame_uart_gcs_group_bin_0156 = frame (4k)
frame_uart_gcs_group_bin_0157 = frame (4k)
frame_uart_gcs_group_bin_0158 = frame (4k)
frame_uart_gcs_group_bin_0160 = frame (4k)
frame_uart_gcs_group_bin_0161 = frame (4k)
frame_uart_gcs_group_bin_0162 = frame (4k)
frame_uart_gcs_group_bin_0163 = frame (4k)
frame_uart_gcs_group_bin_0164 = frame (4k)
frame_uart_gcs_group_bin_0165 = frame (4k)
frame_uart_gcs_group_bin_0166 = frame (4k)
frame_uart_gcs_group_bin_0167 = frame (4k)
frame_uart_gcs_group_bin_0168 = frame (4k)
frame_uart_gcs_group_bin_0169 = frame (4k)
frame_uart_gcs_group_bin_0170 = frame (4k)
frame_uart_gcs_group_bin_0171 = frame (4k)
frame_uart_gcs_group_bin_0172 = frame (4k)
frame_uart_gcs_group_bin_0173 = frame (4k)
frame_uart_gcs_group_bin_0174 = frame (4k)
frame_uart_gcs_group_bin_0175 = frame (4k)
frame_uart_gcs_group_bin_0176 = frame (4k)
frame_uart_gcs_group_bin_0177 = frame (4k)
frame_uart_gcs_group_bin_0178 = frame (4k)
frame_uart_gcs_group_bin_0180 = frame (4k)
frame_uart_gcs_group_bin_0181 = frame (4k)
frame_uart_gcs_group_bin_0182 = frame (4k)
frame_uart_gcs_group_bin_0183 = frame (4k)
frame_uart_gcs_group_bin_0184 = frame (4k)
frame_uart_gcs_group_bin_0185 = frame (4k)
frame_uart_gcs_group_bin_0186 = frame (4k)
frame_uart_gcs_group_bin_0188 = frame (4k)
frame_uart_gcs_group_bin_0189 = frame (4k)
frame_uart_gcs_group_bin_0190 = frame (4k)
frame_uart_gcs_group_bin_0191 = frame (4k)
frame_uart_gcs_group_bin_0192 = frame (4k)
frame_uart_gcs_group_bin_0193 = frame (4k)
frame_uart_gcs_group_bin_0194 = frame (4k)
frame_uart_gcs_group_bin_0196 = frame (4k)
frame_uart_gcs_group_bin_0197 = frame (4k)
frame_uart_gcs_group_bin_0198 = frame (4k)
frame_uart_gcs_group_bin_0199 = frame (4k)
frame_uart_gcs_group_bin_0200 = frame (4k)
frame_uart_gcs_group_bin_0202 = frame (4k)
frame_uart_gcs_group_bin_0203 = frame (4k)
frame_uart_gcs_group_bin_0204 = frame (4k)
frame_uart_gcs_group_bin_0205 = frame (4k)
frame_uart_gcs_group_bin_0206 = frame (4k)
frame_uart_gcs_group_bin_0207 = frame (4k)
frame_uart_gcs_group_bin_0208 = frame (4k)
frame_uart_gcs_group_bin_0209 = frame (4k)
frame_uart_gcs_group_bin_0210 = frame (4k)
frame_uart_gcs_group_bin_0211 = frame (4k)
frame_uart_gcs_group_bin_0212 = frame (4k)
frame_uart_gcs_group_bin_0213 = frame (4k)
frame_uart_gcs_group_bin_0214 = frame (4k)
frame_uart_gcs_group_bin_0215 = frame (4k)
frame_uart_gcs_group_bin_0216 = frame (4k)
frame_uart_gcs_group_bin_0217 = frame (4k)
frame_uart_gcs_group_bin_0218 = frame (4k)
frame_uart_gcs_group_bin_0219 = frame (4k)
frame_uart_gcs_group_bin_0220 = frame (4k)
frame_uart_gcs_group_bin_0221 = frame (4k)
frame_uart_gcs_group_bin_0222 = frame (4k)
frame_uart_gcs_group_bin_0223 = frame (4k)
frame_uart_gcs_group_bin_0224 = frame (4k)
frame_uart_gcs_group_bin_0225 = frame (4k)
frame_uart_gcs_group_bin_0226 = frame (4k)
frame_uart_gcs_group_bin_0227 = frame (4k)
frame_uart_gcs_group_bin_0228 = frame (4k)
frame_uart_gcs_group_bin_0230 = frame (4k)
frame_uart_gcs_group_bin_0231 = frame (4k)
frame_uart_gcs_group_bin_0232 = frame (4k)
frame_uart_gcs_group_bin_0233 = frame (4k)
frame_uart_gcs_group_bin_0234 = frame (4k)
frame_uart_gcs_group_bin_0235 = frame (4k)
frame_uart_gcs_group_bin_0236 = frame (4k)
frame_uart_gcs_group_bin_0237 = frame (4k)
frame_uart_gcs_group_bin_0238 = frame (4k)
frame_uart_gcs_group_bin_0239 = frame (4k)
frame_uart_gcs_group_bin_0240 = frame (4k)
frame_uart_gcs_group_bin_0241 = frame (4k)
frame_uart_gcs_group_bin_0242 = frame (4k)
frame_uart_gcs_group_bin_0243 = frame (4k)
frame_uart_gcs_group_bin_0244 = frame (4k)
frame_uart_gcs_group_bin_0245 = frame (4k, paddr: 0x12c30000)
frame_uart_gcs_group_bin_0246 = frame (4k)
frame_uart_gcs_group_bin_0247 = frame (4k)
frame_uart_gcs_group_bin_0248 = frame (4k)
frame_uart_gcs_group_bin_0249 = frame (4k)
frame_uart_gcs_group_bin_0250 = frame (4k)
frame_uart_gcs_group_bin_0251 = frame (4k)
frame_uart_gcs_group_bin_0252 = frame (4k)
frame_uart_gcs_group_bin_0253 = frame (4k)
frame_uart_gcs_group_bin_0254 = frame (4k)
frame_uart_gcs_group_bin_0255 = frame (4k)
frame_uart_gcs_group_bin_0256 = frame (4k)
frame_uart_gcs_group_bin_0257 = frame (4k)
frame_uart_gcs_group_bin_0258 = frame (4k)
frame_uart_gcs_group_bin_0260 = frame (4k)
frame_uart_gcs_group_bin_0261 = frame (4k)
frame_uart_gcs_group_bin_0262 = frame (4k)
frame_uart_gcs_group_bin_0263 = frame (4k)
frame_uart_gcs_group_bin_0264 = frame (4k)
frame_uart_gcs_group_bin_0265 = frame (4k)
frame_uart_gcs_group_bin_0266 = frame (4k)
frame_uart_gcs_group_bin_0267 = frame (4k)
frame_uart_gcs_group_bin_0269 = frame (4k)
frame_uart_gcs_group_bin_0270 = frame (4k)
frame_uart_gcs_group_bin_0271 = frame (4k)
frame_uart_gcs_group_bin_0272 = frame (4k)
frame_uart_gcs_group_bin_0273 = frame (4k)
frame_uart_gcs_group_bin_0274 = frame (4k)
frame_uart_gcs_group_bin_0275 = frame (4k)
frame_uart_gcs_group_bin_0276 = frame (4k)
frame_uart_gcs_group_bin_0277 = frame (4k)
frame_uart_gcs_group_bin_0278 = frame (4k)
frame_uart_gcs_group_bin_0279 = frame (4k)
frame_uart_gcs_group_bin_0280 = frame (4k)
frame_uart_gcs_group_bin_0281 = frame (4k)
frame_uart_gcs_group_bin_0282 = frame (4k)
frame_uart_gcs_group_bin_0283 = frame (4k)
frame_uart_gcs_group_bin_0284 = frame (4k)
frame_uart_gcs_group_bin_0285 = frame (4k)
frame_uart_gcs_group_bin_0286 = frame (4k)
frame_uart_gcs_group_bin_0287 = frame (4k)
frame_uart_gcs_group_bin_0288 = frame (4k)
frame_uart_gcs_group_bin_0289 = frame (4k)
frame_uart_gcs_group_bin_0290 = frame (4k)
frame_uart_gcs_group_bin_0291 = frame (4k)
frame_uart_gcs_group_bin_0292 = frame (4k)
frame_uart_gcs_group_bin_0293 = frame (4k)
frame_uart_gcs_group_bin_0294 = frame (4k)
frame_uart_gcs_group_bin_0295 = frame (4k)
frame_uart_gcs_group_bin_0296 = frame (4k)
frame_uart_gcs_group_bin_0297 = frame (4k)
frame_uart_gcs_group_bin_0298 = frame (4k)
frame_uart_gcs_group_bin_0299 = frame (4k)
frame_uart_gcs_group_bin_0300 = frame (4k)
frame_uart_gcs_group_bin_0301 = frame (4k)
frame_uart_gcs_group_bin_0302 = frame (4k)
frame_uart_gcs_group_bin_0303 = frame (4k)
frame_uart_gcs_group_bin_0304 = frame (4k)
frame_uart_gcs_group_bin_0305 = frame (4k)
frame_uart_gcs_group_bin_0306 = frame (4k)
frame_uart_gcs_group_bin_0307 = frame (4k)
frame_uart_gcs_group_bin_0308 = frame (4k)
frame_uart_gcs_group_bin_0309 = frame (4k)
frame_uart_gcs_group_bin_0310 = frame (4k)
frame_uart_gcs_group_bin_0311 = frame (4k)
frame_uart_gcs_group_bin_0312 = frame (4k)
frame_uart_gcs_group_bin_0313 = frame (4k)
frame_uart_px4_group_bin_0000 = frame (4k)
frame_uart_px4_group_bin_0001 = frame (4k)
frame_uart_px4_group_bin_0002 = frame (4k)
frame_uart_px4_group_bin_0003 = frame (4k)
frame_uart_px4_group_bin_0004 = frame (4k)
frame_uart_px4_group_bin_0005 = frame (4k)
frame_uart_px4_group_bin_0006 = frame (4k)
frame_uart_px4_group_bin_0007 = frame (4k)
frame_uart_px4_group_bin_0008 = frame (4k)
frame_uart_px4_group_bin_0009 = frame (4k)
frame_uart_px4_group_bin_0010 = frame (4k)
frame_uart_px4_group_bin_0011 = frame (4k)
frame_uart_px4_group_bin_0012 = frame (4k)
frame_uart_px4_group_bin_0013 = frame (4k)
frame_uart_px4_group_bin_0014 = frame (4k)
frame_uart_px4_group_bin_0017 = frame (4k)
frame_uart_px4_group_bin_0018 = frame (4k)
frame_uart_px4_group_bin_0019 = frame (4k)
frame_uart_px4_group_bin_0020 = frame (4k)
frame_uart_px4_group_bin_0021 = frame (4k)
frame_uart_px4_group_bin_0022 = frame (4k)
frame_uart_px4_group_bin_0024 = frame (4k)
frame_uart_px4_group_bin_0025 = frame (4k)
frame_uart_px4_group_bin_0026 = frame (4k)
frame_uart_px4_group_bin_0027 = frame (4k)
frame_uart_px4_group_bin_0028 = frame (4k)
frame_uart_px4_group_bin_0029 = frame (4k)
frame_uart_px4_group_bin_0030 = frame (4k)
frame_uart_px4_group_bin_0031 = frame (4k)
frame_uart_px4_group_bin_0032 = frame (4k)
frame_uart_px4_group_bin_0033 = frame (4k)
frame_uart_px4_group_bin_0034 = frame (4k)
frame_uart_px4_group_bin_0035 = frame (4k)
frame_uart_px4_group_bin_0036 = frame (4k)
frame_uart_px4_group_bin_0037 = frame (4k)
frame_uart_px4_group_bin_0038 = frame (4k)
frame_uart_px4_group_bin_0039 = frame (4k)
frame_uart_px4_group_bin_0040 = frame (4k)
frame_uart_px4_group_bin_0041 = frame (4k)
frame_uart_px4_group_bin_0042 = frame (4k)
frame_uart_px4_group_bin_0043 = frame (4k)
frame_uart_px4_group_bin_0044 = frame (4k)
frame_uart_px4_group_bin_0045 = frame (4k)
frame_uart_px4_group_bin_0046 = frame (4k)
frame_uart_px4_group_bin_0047 = frame (4k)
frame_uart_px4_group_bin_0048 = frame (4k)
frame_uart_px4_group_bin_0049 = frame (4k)
frame_uart_px4_group_bin_0050 = frame (4k)
frame_uart_px4_group_bin_0051 = frame (4k)
frame_uart_px4_group_bin_0052 = frame (4k)
frame_uart_px4_group_bin_0053 = frame (4k)
frame_uart_px4_group_bin_0054 = frame (4k)
frame_uart_px4_group_bin_0055 = frame (4k)
frame_uart_px4_group_bin_0057 = frame (4k)
frame_uart_px4_group_bin_0059 = frame (4k)
frame_uart_px4_group_bin_0060 = frame (4k)
frame_uart_px4_group_bin_0061 = frame (4k)
frame_uart_px4_group_bin_0062 = frame (4k)
frame_uart_px4_group_bin_0063 = frame (4k)
frame_uart_px4_group_bin_0064 = frame (4k)
frame_uart_px4_group_bin_0065 = frame (4k)
frame_uart_px4_group_bin_0066 = frame (4k)
frame_uart_px4_group_bin_0067 = frame (4k)
frame_uart_px4_group_bin_0068 = frame (4k)
frame_uart_px4_group_bin_0069 = frame (4k)
frame_uart_px4_group_bin_0070 = frame (4k)
frame_uart_px4_group_bin_0071 = frame (4k)
frame_uart_px4_group_bin_0072 = frame (4k)
frame_uart_px4_group_bin_0073 = frame (4k)
frame_uart_px4_group_bin_0074 = frame (4k)
frame_uart_px4_group_bin_0075 = frame (4k)
frame_uart_px4_group_bin_0076 = frame (4k)
frame_uart_px4_group_bin_0077 = frame (4k)
frame_uart_px4_group_bin_0078 = frame (4k)
frame_uart_px4_group_bin_0079 = frame (4k)
frame_uart_px4_group_bin_0080 = frame (4k)
frame_uart_px4_group_bin_0081 = frame (4k)
frame_uart_px4_group_bin_0082 = frame (4k)
frame_uart_px4_group_bin_0083 = frame (4k)
frame_uart_px4_group_bin_0084 = frame (4k)
frame_uart_px4_group_bin_0085 = frame (4k)
frame_uart_px4_group_bin_0086 = frame (4k)
frame_uart_px4_group_bin_0087 = frame (4k)
frame_uart_px4_group_bin_0088 = frame (4k)
frame_uart_px4_group_bin_0089 = frame (4k)
frame_uart_px4_group_bin_0090 = frame (4k)
frame_uart_px4_group_bin_0091 = frame (4k)
frame_uart_px4_group_bin_0092 = frame (4k)
frame_uart_px4_group_bin_0093 = frame (4k)
frame_uart_px4_group_bin_0094 = frame (4k)
frame_uart_px4_group_bin_0095 = frame (4k)
frame_uart_px4_group_bin_0096 = frame (4k)
frame_uart_px4_group_bin_0097 = frame (4k)
frame_uart_px4_group_bin_0098 = frame (4k)
frame_uart_px4_group_bin_0099 = frame (4k)
frame_uart_px4_group_bin_0100 = frame (4k)
frame_uart_px4_group_bin_0101 = frame (4k)
frame_uart_px4_group_bin_0102 = frame (4k)
frame_uart_px4_group_bin_0104 = frame (4k)
frame_uart_px4_group_bin_0105 = frame (4k)
frame_uart_px4_group_bin_0106 = frame (4k)
frame_uart_px4_group_bin_0107 = frame (4k)
frame_uart_px4_group_bin_0108 = frame (4k)
frame_uart_px4_group_bin_0109 = frame (4k)
frame_uart_px4_group_bin_0110 = frame (4k)
frame_uart_px4_group_bin_0111 = frame (4k)
frame_uart_px4_group_bin_0112 = frame (4k)
frame_uart_px4_group_bin_0113 = frame (4k)
frame_uart_px4_group_bin_0114 = frame (4k)
frame_uart_px4_group_bin_0115 = frame (4k)
frame_uart_px4_group_bin_0116 = frame (4k)
frame_uart_px4_group_bin_0117 = frame (4k)
frame_uart_px4_group_bin_0118 = frame (4k)
frame_uart_px4_group_bin_0119 = frame (4k)
frame_uart_px4_group_bin_0120 = frame (4k)
frame_uart_px4_group_bin_0121 = frame (4k)
frame_uart_px4_group_bin_0122 = frame (4k)
frame_uart_px4_group_bin_0123 = frame (4k)
frame_uart_px4_group_bin_0124 = frame (4k)
frame_uart_px4_group_bin_0125 = frame (4k)
frame_uart_px4_group_bin_0126 = frame (4k)
frame_uart_px4_group_bin_0128 = frame (4k)
frame_uart_px4_group_bin_0129 = frame (4k)
frame_uart_px4_group_bin_0130 = frame (4k)
frame_uart_px4_group_bin_0131 = frame (4k)
frame_uart_px4_group_bin_0132 = frame (4k)
frame_uart_px4_group_bin_0133 = frame (4k)
frame_uart_px4_group_bin_0134 = frame (4k)
frame_uart_px4_group_bin_0135 = frame (4k)
frame_uart_px4_group_bin_0136 = frame (4k)
frame_uart_px4_group_bin_0137 = frame (4k)
frame_uart_px4_group_bin_0138 = frame (4k)
frame_uart_px4_group_bin_0139 = frame (4k)
frame_uart_px4_group_bin_0140 = frame (4k)
frame_uart_px4_group_bin_0141 = frame (4k)
frame_uart_px4_group_bin_0142 = frame (4k)
frame_uart_px4_group_bin_0143 = frame (4k)
frame_uart_px4_group_bin_0145 = frame (4k)
frame_uart_px4_group_bin_0146 = frame (4k)
frame_uart_px4_group_bin_0147 = frame (4k)
frame_uart_px4_group_bin_0148 = frame (4k)
frame_uart_px4_group_bin_0149 = frame (4k)
frame_uart_px4_group_bin_0150 = frame (4k)
frame_uart_px4_group_bin_0151 = frame (4k)
frame_uart_px4_group_bin_0152 = frame (4k)
frame_uart_px4_group_bin_0153 = frame (4k)
frame_uart_px4_group_bin_0154 = frame (4k)
frame_uart_px4_group_bin_0155 = frame (4k)
frame_uart_px4_group_bin_0156 = frame (4k)
frame_uart_px4_group_bin_0157 = frame (4k)
frame_uart_px4_group_bin_0158 = frame (4k)
frame_uart_px4_group_bin_0160 = frame (4k)
frame_uart_px4_group_bin_0161 = frame (4k)
frame_uart_px4_group_bin_0162 = frame (4k)
frame_uart_px4_group_bin_0163 = frame (4k)
frame_uart_px4_group_bin_0164 = frame (4k)
frame_uart_px4_group_bin_0165 = frame (4k)
frame_uart_px4_group_bin_0166 = frame (4k)
frame_uart_px4_group_bin_0167 = frame (4k)
frame_uart_px4_group_bin_0168 = frame (4k)
frame_uart_px4_group_bin_0169 = frame (4k)
frame_uart_px4_group_bin_0171 = frame (4k)
frame_uart_px4_group_bin_0172 = frame (4k)
frame_uart_px4_group_bin_0173 = frame (4k)
frame_uart_px4_group_bin_0174 = frame (4k)
frame_uart_px4_group_bin_0175 = frame (4k)
frame_uart_px4_group_bin_0176 = frame (4k)
frame_uart_px4_group_bin_0177 = frame (4k)
frame_uart_px4_group_bin_0178 = frame (4k)
frame_uart_px4_group_bin_0180 = frame (4k)
frame_uart_px4_group_bin_0181 = frame (4k)
frame_uart_px4_group_bin_0182 = frame (4k)
frame_uart_px4_group_bin_0183 = frame (4k)
frame_uart_px4_group_bin_0184 = frame (4k)
frame_uart_px4_group_bin_0185 = frame (4k)
frame_uart_px4_group_bin_0186 = frame (4k)
frame_uart_px4_group_bin_0188 = frame (4k)
frame_uart_px4_group_bin_0189 = frame (4k)
frame_uart_px4_group_bin_0190 = frame (4k)
frame_uart_px4_group_bin_0191 = frame (4k)
frame_uart_px4_group_bin_0192 = frame (4k)
frame_uart_px4_group_bin_0193 = frame (4k)
frame_uart_px4_group_bin_0194 = frame (4k)
frame_uart_px4_group_bin_0196 = frame (4k)
frame_uart_px4_group_bin_0197 = frame (4k)
frame_uart_px4_group_bin_0198 = frame (4k)
frame_uart_px4_group_bin_0199 = frame (4k)
frame_uart_px4_group_bin_0200 = frame (4k)
frame_uart_px4_group_bin_0202 = frame (4k)
frame_uart_px4_group_bin_0203 = frame (4k)
frame_uart_px4_group_bin_0204 = frame (4k)
frame_uart_px4_group_bin_0205 = frame (4k)
frame_uart_px4_group_bin_0206 = frame (4k)
frame_uart_px4_group_bin_0207 = frame (4k)
frame_uart_px4_group_bin_0208 = frame (4k)
frame_uart_px4_group_bin_0209 = frame (4k)
frame_uart_px4_group_bin_0210 = frame (4k)
frame_uart_px4_group_bin_0211 = frame (4k)
frame_uart_px4_group_bin_0212 = frame (4k)
frame_uart_px4_group_bin_0213 = frame (4k)
frame_uart_px4_group_bin_0214 = frame (4k)
frame_uart_px4_group_bin_0215 = frame (4k)
frame_uart_px4_group_bin_0216 = frame (4k)
frame_uart_px4_group_bin_0217 = frame (4k)
frame_uart_px4_group_bin_0218 = frame (4k)
frame_uart_px4_group_bin_0219 = frame (4k)
frame_uart_px4_group_bin_0220 = frame (4k)
frame_uart_px4_group_bin_0221 = frame (4k)
frame_uart_px4_group_bin_0222 = frame (4k)
frame_uart_px4_group_bin_0223 = frame (4k)
frame_uart_px4_group_bin_0224 = frame (4k)
frame_uart_px4_group_bin_0225 = frame (4k)
frame_uart_px4_group_bin_0226 = frame (4k)
frame_uart_px4_group_bin_0227 = frame (4k)
frame_uart_px4_group_bin_0228 = frame (4k)
frame_uart_px4_group_bin_0230 = frame (4k)
frame_uart_px4_group_bin_0231 = frame (4k)
frame_uart_px4_group_bin_0232 = frame (4k)
frame_uart_px4_group_bin_0233 = frame (4k)
frame_uart_px4_group_bin_0234 = frame (4k)
frame_uart_px4_group_bin_0235 = frame (4k)
frame_uart_px4_group_bin_0236 = frame (4k)
frame_uart_px4_group_bin_0237 = frame (4k)
frame_uart_px4_group_bin_0238 = frame (4k)
frame_uart_px4_group_bin_0239 = frame (4k)
frame_uart_px4_group_bin_0240 = frame (4k)
frame_uart_px4_group_bin_0241 = frame (4k)
frame_uart_px4_group_bin_0242 = frame (4k)
frame_uart_px4_group_bin_0243 = frame (4k)
frame_uart_px4_group_bin_0244 = frame (4k)
frame_uart_px4_group_bin_0245 = frame (4k, paddr: 0x12c10000)
frame_uart_px4_group_bin_0246 = frame (4k)
frame_uart_px4_group_bin_0247 = frame (4k)
frame_uart_px4_group_bin_0248 = frame (4k)
frame_uart_px4_group_bin_0249 = frame (4k)
frame_uart_px4_group_bin_0250 = frame (4k)
frame_uart_px4_group_bin_0251 = frame (4k)
frame_uart_px4_group_bin_0252 = frame (4k)
frame_uart_px4_group_bin_0253 = frame (4k)
frame_uart_px4_group_bin_0254 = frame (4k)
frame_uart_px4_group_bin_0255 = frame (4k)
frame_uart_px4_group_bin_0256 = frame (4k)
frame_uart_px4_group_bin_0257 = frame (4k)
frame_uart_px4_group_bin_0258 = frame (4k)
frame_uart_px4_group_bin_0260 = frame (4k)
frame_uart_px4_group_bin_0261 = frame (4k)
frame_uart_px4_group_bin_0262 = frame (4k)
frame_uart_px4_group_bin_0263 = frame (4k)
frame_uart_px4_group_bin_0264 = frame (4k)
frame_uart_px4_group_bin_0265 = frame (4k)
frame_uart_px4_group_bin_0266 = frame (4k)
frame_uart_px4_group_bin_0267 = frame (4k)
frame_uart_px4_group_bin_0269 = frame (4k)
frame_uart_px4_group_bin_0270 = frame (4k)
frame_uart_px4_group_bin_0271 = frame (4k)
frame_uart_px4_group_bin_0272 = frame (4k)
frame_uart_px4_group_bin_0273 = frame (4k)
frame_uart_px4_group_bin_0274 = frame (4k)
frame_uart_px4_group_bin_0275 = frame (4k)
frame_uart_px4_group_bin_0276 = frame (4k)
frame_uart_px4_group_bin_0277 = frame (4k)
frame_uart_px4_group_bin_0278 = frame (4k)
frame_uart_px4_group_bin_0279 = frame (4k)
frame_uart_px4_group_bin_0280 = frame (4k)
frame_uart_px4_group_bin_0281 = frame (4k)
frame_uart_px4_group_bin_0282 = frame (4k)
frame_uart_px4_group_bin_0283 = frame (4k)
frame_uart_px4_group_bin_0284 = frame (4k)
frame_uart_px4_group_bin_0285 = frame (4k)
frame_uart_px4_group_bin_0286 = frame (4k)
frame_uart_px4_group_bin_0287 = frame (4k)
frame_uart_px4_group_bin_0288 = frame (4k)
frame_uart_px4_group_bin_0289 = frame (4k)
frame_uart_px4_group_bin_0290 = frame (4k)
frame_uart_px4_group_bin_0291 = frame (4k)
frame_uart_px4_group_bin_0292 = frame (4k)
frame_uart_px4_group_bin_0293 = frame (4k)
frame_uart_px4_group_bin_0294 = frame (4k)
frame_uart_px4_group_bin_0295 = frame (4k)
frame_uart_px4_group_bin_0296 = frame (4k)
frame_uart_px4_group_bin_0297 = frame (4k)
frame_uart_px4_group_bin_0298 = frame (4k)
frame_uart_px4_group_bin_0299 = frame (4k)
frame_uart_px4_group_bin_0300 = frame (4k)
frame_uart_px4_group_bin_0301 = frame (4k)
frame_uart_px4_group_bin_0302 = frame (4k)
frame_uart_px4_group_bin_0303 = frame (4k)
frame_uart_px4_group_bin_0304 = frame (4k)
frame_uart_px4_group_bin_0305 = frame (4k)
frame_uart_px4_group_bin_0306 = frame (4k)
frame_uart_px4_group_bin_0307 = frame (4k)
frame_uart_px4_group_bin_0308 = frame (4k)
frame_uart_px4_group_bin_0309 = frame (4k)
frame_uart_px4_group_bin_0310 = frame (4k)
frame_uart_px4_group_bin_0311 = frame (4k)
frame_uart_px4_group_bin_0312 = frame (4k)
frame_uart_px4_group_bin_0313 = frame (4k)
frame_vm_group_bin_0000 = frame (4k)
frame_vm_group_bin_0001 = frame (4k)
frame_vm_group_bin_0002 = frame (4k)
frame_vm_group_bin_0003 = frame (4k)
frame_vm_group_bin_0004 = frame (4k)
frame_vm_group_bin_0005 = frame (4k)
frame_vm_group_bin_0006 = frame (4k)
frame_vm_group_bin_0007 = frame (4k)
frame_vm_group_bin_0008 = frame (4k)
frame_vm_group_bin_0009 = frame (4k)
frame_vm_group_bin_0010 = frame (4k)
frame_vm_group_bin_0011 = frame (4k)
frame_vm_group_bin_0012 = frame (4k)
frame_vm_group_bin_0013 = frame (4k)
frame_vm_group_bin_0014 = frame (4k)
frame_vm_group_bin_0015 = frame (4k)
frame_vm_group_bin_0016 = frame (4k)
frame_vm_group_bin_0017 = frame (4k)
frame_vm_group_bin_0018 = frame (4k)
frame_vm_group_bin_0019 = frame (4k)
frame_vm_group_bin_0020 = frame (4k)
frame_vm_group_bin_0021 = frame (4k)
frame_vm_group_bin_0022 = frame (4k)
frame_vm_group_bin_0023 = frame (4k)
frame_vm_group_bin_0024 = frame (4k)
frame_vm_group_bin_0025 = frame (4k)
frame_vm_group_bin_0026 = frame (4k)
frame_vm_group_bin_0027 = frame (4k)
frame_vm_group_bin_0028 = frame (4k)
frame_vm_group_bin_0029 = frame (4k)
frame_vm_group_bin_0030 = frame (4k)
frame_vm_group_bin_0031 = frame (4k)
frame_vm_group_bin_0032 = frame (4k)
frame_vm_group_bin_0033 = frame (4k)
frame_vm_group_bin_0034 = frame (4k)
frame_vm_group_bin_0035 = frame (4k)
frame_vm_group_bin_0036 = frame (4k)
frame_vm_group_bin_0037 = frame (4k)
frame_vm_group_bin_0038 = frame (4k)
frame_vm_group_bin_0039 = frame (4k)
frame_vm_group_bin_0040 = frame (4k)
frame_vm_group_bin_0041 = frame (4k)
frame_vm_group_bin_0042 = frame (4k)
frame_vm_group_bin_0043 = frame (4k)
frame_vm_group_bin_0044 = frame (4k)
frame_vm_group_bin_0045 = frame (4k)
frame_vm_group_bin_0046 = frame (4k)
frame_vm_group_bin_0047 = frame (4k)
frame_vm_group_bin_0048 = frame (4k)
frame_vm_group_bin_0049 = frame (4k)
frame_vm_group_bin_0050 = frame (4k)
frame_vm_group_bin_0051 = frame (4k)
frame_vm_group_bin_0052 = frame (4k)
frame_vm_group_bin_0053 = frame (4k)
frame_vm_group_bin_0054 = frame (4k)
frame_vm_group_bin_0055 = frame (4k)
frame_vm_group_bin_0056 = frame (4k)
frame_vm_group_bin_0057 = frame (4k)
frame_vm_group_bin_0058 = frame (4k)
frame_vm_group_bin_0059 = frame (4k)
frame_vm_group_bin_0060 = frame (4k)
frame_vm_group_bin_0061 = frame (4k)
frame_vm_group_bin_0062 = frame (4k)
frame_vm_group_bin_0063 = frame (4k)
frame_vm_group_bin_0064 = frame (4k)
frame_vm_group_bin_0065 = frame (4k)
frame_vm_group_bin_0066 = frame (4k)
frame_vm_group_bin_0067 = frame (4k)
frame_vm_group_bin_0068 = frame (4k)
frame_vm_group_bin_0069 = frame (4k)
frame_vm_group_bin_0070 = frame (4k)
frame_vm_group_bin_0071 = frame (4k)
frame_vm_group_bin_0072 = frame (4k)
frame_vm_group_bin_0073 = frame (4k)
frame_vm_group_bin_0074 = frame (4k)
frame_vm_group_bin_0075 = frame (4k)
frame_vm_group_bin_0076 = frame (4k)
frame_vm_group_bin_0077 = frame (4k)
frame_vm_group_bin_0078 = frame (4k)
frame_vm_group_bin_0079 = frame (4k)
frame_vm_group_bin_0080 = frame (4k)
frame_vm_group_bin_0081 = frame (4k)
frame_vm_group_bin_0082 = frame (4k)
frame_vm_group_bin_0083 = frame (4k)
frame_vm_group_bin_0084 = frame (4k)
frame_vm_group_bin_0085 = frame (4k)
frame_vm_group_bin_0086 = frame (4k)
frame_vm_group_bin_0087 = frame (4k)
frame_vm_group_bin_0088 = frame (4k)
frame_vm_group_bin_0089 = frame (4k)
frame_vm_group_bin_0090 = frame (4k)
frame_vm_group_bin_0091 = frame (4k)
frame_vm_group_bin_0092 = frame (4k)
frame_vm_group_bin_0093 = frame (4k)
frame_vm_group_bin_0094 = frame (4k)
frame_vm_group_bin_0095 = frame (4k)
frame_vm_group_bin_0096 = frame (4k)
frame_vm_group_bin_0097 = frame (4k)
frame_vm_group_bin_0098 = frame (4k)
frame_vm_group_bin_0099 = frame (4k)
frame_vm_group_bin_0100 = frame (4k)
frame_vm_group_bin_0101 = frame (4k)
frame_vm_group_bin_0102 = frame (4k)
frame_vm_group_bin_0103 = frame (4k)
frame_vm_group_bin_0104 = frame (4k)
frame_vm_group_bin_0105 = frame (4k)
frame_vm_group_bin_0106 = frame (4k)
frame_vm_group_bin_0107 = frame (4k)
frame_vm_group_bin_0108 = frame (4k)
frame_vm_group_bin_0109 = frame (4k)
frame_vm_group_bin_0110 = frame (4k)
frame_vm_group_bin_0111 = frame (4k)
frame_vm_group_bin_0112 = frame (4k)
frame_vm_group_bin_0113 = frame (4k)
frame_vm_group_bin_0114 = frame (4k)
frame_vm_group_bin_0115 = frame (4k)
frame_vm_group_bin_0116 = frame (4k)
frame_vm_group_bin_0117 = frame (4k)
frame_vm_group_bin_0118 = frame (4k)
frame_vm_group_bin_0119 = frame (4k)
frame_vm_group_bin_0120 = frame (4k)
frame_vm_group_bin_0121 = frame (4k)
frame_vm_group_bin_0122 = frame (4k)
frame_vm_group_bin_0123 = frame (4k)
frame_vm_group_bin_0124 = frame (4k)
frame_vm_group_bin_0125 = frame (4k)
frame_vm_group_bin_0126 = frame (4k)
frame_vm_group_bin_0127 = frame (4k)
frame_vm_group_bin_0128 = frame (4k)
frame_vm_group_bin_0129 = frame (4k)
frame_vm_group_bin_0130 = frame (4k)
frame_vm_group_bin_0131 = frame (4k)
frame_vm_group_bin_0132 = frame (4k)
frame_vm_group_bin_0133 = frame (4k)
frame_vm_group_bin_0134 = frame (4k)
frame_vm_group_bin_0135 = frame (4k)
frame_vm_group_bin_0136 = frame (4k)
frame_vm_group_bin_0137 = frame (4k)
frame_vm_group_bin_0138 = frame (4k)
frame_vm_group_bin_0139 = frame (4k)
frame_vm_group_bin_0140 = frame (4k)
frame_vm_group_bin_0141 = frame (4k)
frame_vm_group_bin_0142 = frame (4k)
frame_vm_group_bin_0143 = frame (4k)
frame_vm_group_bin_0144 = frame (4k)
frame_vm_group_bin_0145 = frame (4k)
frame_vm_group_bin_0146 = frame (4k)
frame_vm_group_bin_0147 = frame (4k)
frame_vm_group_bin_0148 = frame (4k)
frame_vm_group_bin_0149 = frame (4k)
frame_vm_group_bin_0150 = frame (4k)
frame_vm_group_bin_0151 = frame (4k)
frame_vm_group_bin_0152 = frame (4k)
frame_vm_group_bin_0153 = frame (4k)
frame_vm_group_bin_0154 = frame (4k)
frame_vm_group_bin_0155 = frame (4k)
frame_vm_group_bin_0156 = frame (4k)
frame_vm_group_bin_0157 = frame (4k)
frame_vm_group_bin_0158 = frame (4k)
frame_vm_group_bin_0159 = frame (4k)
frame_vm_group_bin_0160 = frame (4k)
frame_vm_group_bin_0161 = frame (4k)
frame_vm_group_bin_0162 = frame (4k)
frame_vm_group_bin_0163 = frame (4k)
frame_vm_group_bin_0164 = frame (4k)
frame_vm_group_bin_0165 = frame (4k)
frame_vm_group_bin_0166 = frame (4k)
frame_vm_group_bin_0167 = frame (4k)
frame_vm_group_bin_0168 = frame (4k)
frame_vm_group_bin_0169 = frame (4k)
frame_vm_group_bin_0170 = frame (4k)
frame_vm_group_bin_0171 = frame (4k)
frame_vm_group_bin_0172 = frame (4k)
frame_vm_group_bin_0173 = frame (4k)
frame_vm_group_bin_0174 = frame (4k)
frame_vm_group_bin_0175 = frame (4k)
frame_vm_group_bin_0176 = frame (4k)
frame_vm_group_bin_0177 = frame (4k)
frame_vm_group_bin_0178 = frame (4k)
frame_vm_group_bin_0179 = frame (4k)
frame_vm_group_bin_0180 = frame (4k)
frame_vm_group_bin_0181 = frame (4k)
frame_vm_group_bin_0182 = frame (4k)
frame_vm_group_bin_0183 = frame (4k)
frame_vm_group_bin_0184 = frame (4k)
frame_vm_group_bin_0185 = frame (4k)
frame_vm_group_bin_0186 = frame (4k)
frame_vm_group_bin_0187 = frame (4k)
frame_vm_group_bin_0188 = frame (4k)
frame_vm_group_bin_0189 = frame (4k)
frame_vm_group_bin_0190 = frame (4k)
frame_vm_group_bin_0191 = frame (4k)
frame_vm_group_bin_0192 = frame (4k)
frame_vm_group_bin_0193 = frame (4k)
frame_vm_group_bin_0194 = frame (4k)
frame_vm_group_bin_0195 = frame (4k)
frame_vm_group_bin_0196 = frame (4k)
frame_vm_group_bin_0197 = frame (4k)
frame_vm_group_bin_0198 = frame (4k)
frame_vm_group_bin_0199 = frame (4k)
frame_vm_group_bin_0200 = frame (4k)
frame_vm_group_bin_0201 = frame (4k)
frame_vm_group_bin_0202 = frame (4k)
frame_vm_group_bin_0203 = frame (4k)
frame_vm_group_bin_0204 = frame (4k)
frame_vm_group_bin_0205 = frame (4k)
frame_vm_group_bin_0206 = frame (4k)
frame_vm_group_bin_0207 = frame (4k)
frame_vm_group_bin_0208 = frame (4k)
frame_vm_group_bin_0209 = frame (4k)
frame_vm_group_bin_0210 = frame (4k)
frame_vm_group_bin_0211 = frame (4k)
frame_vm_group_bin_0212 = frame (4k)
frame_vm_group_bin_0213 = frame (4k)
frame_vm_group_bin_0214 = frame (4k)
frame_vm_group_bin_0215 = frame (4k)
frame_vm_group_bin_0216 = frame (4k)
frame_vm_group_bin_0217 = frame (4k)
frame_vm_group_bin_0218 = frame (4k)
frame_vm_group_bin_0219 = frame (4k)
frame_vm_group_bin_0220 = frame (4k)
frame_vm_group_bin_0221 = frame (4k)
frame_vm_group_bin_0222 = frame (4k)
frame_vm_group_bin_0223 = frame (4k)
frame_vm_group_bin_0224 = frame (4k)
frame_vm_group_bin_0225 = frame (4k)
frame_vm_group_bin_0226 = frame (4k)
frame_vm_group_bin_0227 = frame (4k)
frame_vm_group_bin_0228 = frame (4k)
frame_vm_group_bin_0229 = frame (4k)
frame_vm_group_bin_0230 = frame (4k)
frame_vm_group_bin_0231 = frame (4k)
frame_vm_group_bin_0232 = frame (4k)
frame_vm_group_bin_0233 = frame (4k)
frame_vm_group_bin_0234 = frame (4k)
frame_vm_group_bin_0235 = frame (4k)
frame_vm_group_bin_0236 = frame (4k)
frame_vm_group_bin_0237 = frame (4k)
frame_vm_group_bin_0238 = frame (4k)
frame_vm_group_bin_0239 = frame (4k)
frame_vm_group_bin_0240 = frame (4k)
frame_vm_group_bin_0241 = frame (4k)
frame_vm_group_bin_0242 = frame (4k)
frame_vm_group_bin_0243 = frame (4k)
frame_vm_group_bin_0244 = frame (4k)
frame_vm_group_bin_0245 = frame (4k)
frame_vm_group_bin_0246 = frame (4k)
frame_vm_group_bin_0247 = frame (4k)
frame_vm_group_bin_0248 = frame (4k)
frame_vm_group_bin_0249 = frame (4k)
frame_vm_group_bin_0250 = frame (4k)
frame_vm_group_bin_0251 = frame (4k)
frame_vm_group_bin_0252 = frame (4k)
frame_vm_group_bin_0253 = frame (4k)
frame_vm_group_bin_0254 = frame (4k)
frame_vm_group_bin_0255 = frame (4k)
frame_vm_group_bin_0256 = frame (4k)
frame_vm_group_bin_0257 = frame (4k)
frame_vm_group_bin_0258 = frame (4k)
frame_vm_group_bin_0259 = frame (4k)
frame_vm_group_bin_0260 = frame (4k)
frame_vm_group_bin_0261 = frame (4k)
frame_vm_group_bin_0262 = frame (4k)
frame_vm_group_bin_0263 = frame (4k)
frame_vm_group_bin_0264 = frame (4k)
frame_vm_group_bin_0265 = frame (4k)
frame_vm_group_bin_0266 = frame (4k)
frame_vm_group_bin_0267 = frame (4k)
frame_vm_group_bin_0268 = frame (4k)
frame_vm_group_bin_0269 = frame (4k)
frame_vm_group_bin_0270 = frame (4k)
frame_vm_group_bin_0271 = frame (4k)
frame_vm_group_bin_0272 = frame (4k)
frame_vm_group_bin_0273 = frame (4k)
frame_vm_group_bin_0274 = frame (4k)
frame_vm_group_bin_0275 = frame (4k)
frame_vm_group_bin_0276 = frame (4k)
frame_vm_group_bin_0277 = frame (4k)
frame_vm_group_bin_0278 = frame (4k)
frame_vm_group_bin_0279 = frame (4k)
frame_vm_group_bin_0280 = frame (4k)
frame_vm_group_bin_0281 = frame (4k)
frame_vm_group_bin_0282 = frame (4k)
frame_vm_group_bin_0283 = frame (4k)
frame_vm_group_bin_0284 = frame (4k)
frame_vm_group_bin_0285 = frame (4k)
frame_vm_group_bin_0286 = frame (4k)
frame_vm_group_bin_0287 = frame (4k)
frame_vm_group_bin_0288 = frame (4k)
frame_vm_group_bin_0289 = frame (4k)
frame_vm_group_bin_0290 = frame (4k)
frame_vm_group_bin_0291 = frame (4k)
frame_vm_group_bin_0292 = frame (4k)
frame_vm_group_bin_0293 = frame (4k)
frame_vm_group_bin_0294 = frame (4k)
frame_vm_group_bin_0295 = frame (4k)
frame_vm_group_bin_0296 = frame (4k)
frame_vm_group_bin_0297 = frame (4k)
frame_vm_group_bin_0298 = frame (4k)
frame_vm_group_bin_0299 = frame (4k)
frame_vm_group_bin_0300 = frame (4k)
frame_vm_group_bin_0301 = frame (4k)
frame_vm_group_bin_0302 = frame (4k)
frame_vm_group_bin_0303 = frame (4k)
frame_vm_group_bin_0304 = frame (4k)
frame_vm_group_bin_0305 = frame (4k)
frame_vm_group_bin_0306 = frame (4k)
frame_vm_group_bin_0307 = frame (4k)
frame_vm_group_bin_0308 = frame (4k)
frame_vm_group_bin_0309 = frame (4k)
frame_vm_group_bin_0310 = frame (4k)
frame_vm_group_bin_0311 = frame (4k)
frame_vm_group_bin_0312 = frame (4k)
frame_vm_group_bin_0313 = frame (4k)
frame_vm_group_bin_0314 = frame (4k)
frame_vm_group_bin_0315 = frame (4k)
frame_vm_group_bin_0316 = frame (4k)
frame_vm_group_bin_0317 = frame (4k)
frame_vm_group_bin_0318 = frame (4k)
frame_vm_group_bin_0319 = frame (4k)
frame_vm_group_bin_0320 = frame (4k)
frame_vm_group_bin_0321 = frame (4k)
frame_vm_group_bin_0322 = frame (4k)
frame_vm_group_bin_0323 = frame (4k)
frame_vm_group_bin_0324 = frame (4k)
frame_vm_group_bin_0325 = frame (4k)
frame_vm_group_bin_0326 = frame (4k)
frame_vm_group_bin_0327 = frame (4k)
frame_vm_group_bin_0328 = frame (4k)
frame_vm_group_bin_0329 = frame (4k)
frame_vm_group_bin_0330 = frame (4k)
frame_vm_group_bin_0331 = frame (4k)
frame_vm_group_bin_0332 = frame (4k)
frame_vm_group_bin_0333 = frame (4k)
frame_vm_group_bin_0334 = frame (4k)
frame_vm_group_bin_0335 = frame (4k)
frame_vm_group_bin_0336 = frame (4k)
frame_vm_group_bin_0337 = frame (4k)
frame_vm_group_bin_0338 = frame (4k)
frame_vm_group_bin_0339 = frame (4k)
frame_vm_group_bin_0340 = frame (4k)
frame_vm_group_bin_0341 = frame (4k)
frame_vm_group_bin_0342 = frame (4k)
frame_vm_group_bin_0343 = frame (4k)
frame_vm_group_bin_0344 = frame (4k)
frame_vm_group_bin_0345 = frame (4k)
frame_vm_group_bin_0346 = frame (4k)
frame_vm_group_bin_0347 = frame (4k)
frame_vm_group_bin_0348 = frame (4k)
frame_vm_group_bin_0349 = frame (4k)
frame_vm_group_bin_0350 = frame (4k)
frame_vm_group_bin_0351 = frame (4k)
frame_vm_group_bin_0352 = frame (4k)
frame_vm_group_bin_0353 = frame (4k)
frame_vm_group_bin_0354 = frame (4k)
frame_vm_group_bin_0355 = frame (4k)
frame_vm_group_bin_0356 = frame (4k)
frame_vm_group_bin_0357 = frame (4k)
frame_vm_group_bin_0358 = frame (4k)
frame_vm_group_bin_0359 = frame (4k)
frame_vm_group_bin_0360 = frame (4k)
frame_vm_group_bin_0361 = frame (4k)
frame_vm_group_bin_0362 = frame (4k)
frame_vm_group_bin_0363 = frame (4k)
frame_vm_group_bin_0364 = frame (4k)
frame_vm_group_bin_0365 = frame (4k)
frame_vm_group_bin_0366 = frame (4k)
frame_vm_group_bin_0367 = frame (4k)
frame_vm_group_bin_0368 = frame (4k)
frame_vm_group_bin_0369 = frame (4k)
frame_vm_group_bin_0370 = frame (4k)
frame_vm_group_bin_0371 = frame (4k)
frame_vm_group_bin_0372 = frame (4k)
frame_vm_group_bin_0373 = frame (4k)
frame_vm_group_bin_0374 = frame (4k)
frame_vm_group_bin_0375 = frame (4k)
frame_vm_group_bin_0376 = frame (4k)
frame_vm_group_bin_0377 = frame (4k)
frame_vm_group_bin_0378 = frame (4k)
frame_vm_group_bin_0379 = frame (4k)
frame_vm_group_bin_0380 = frame (4k)
frame_vm_group_bin_0381 = frame (4k)
frame_vm_group_bin_0382 = frame (4k)
frame_vm_group_bin_0383 = frame (4k)
frame_vm_group_bin_0384 = frame (4k)
frame_vm_group_bin_0385 = frame (4k)
frame_vm_group_bin_0386 = frame (4k)
frame_vm_group_bin_0387 = frame (4k)
frame_vm_group_bin_0388 = frame (4k)
frame_vm_group_bin_0389 = frame (4k)
frame_vm_group_bin_0390 = frame (4k)
frame_vm_group_bin_0391 = frame (4k)
frame_vm_group_bin_0392 = frame (4k)
frame_vm_group_bin_0393 = frame (4k)
frame_vm_group_bin_0394 = frame (4k)
frame_vm_group_bin_0395 = frame (4k)
frame_vm_group_bin_0396 = frame (4k)
frame_vm_group_bin_0397 = frame (4k)
frame_vm_group_bin_0398 = frame (4k)
frame_vm_group_bin_0399 = frame (4k)
frame_vm_group_bin_0400 = frame (4k)
frame_vm_group_bin_0401 = frame (4k)
frame_vm_group_bin_0402 = frame (4k)
frame_vm_group_bin_0403 = frame (4k)
frame_vm_group_bin_0404 = frame (4k)
frame_vm_group_bin_0405 = frame (4k)
frame_vm_group_bin_0406 = frame (4k)
frame_vm_group_bin_0407 = frame (4k)
frame_vm_group_bin_0408 = frame (4k)
frame_vm_group_bin_0409 = frame (4k)
frame_vm_group_bin_0410 = frame (4k)
frame_vm_group_bin_0411 = frame (4k)
frame_vm_group_bin_0412 = frame (4k)
frame_vm_group_bin_0413 = frame (4k)
frame_vm_group_bin_0414 = frame (4k)
frame_vm_group_bin_0415 = frame (4k)
frame_vm_group_bin_0416 = frame (4k)
frame_vm_group_bin_0417 = frame (4k)
frame_vm_group_bin_0418 = frame (4k)
frame_vm_group_bin_0419 = frame (4k)
frame_vm_group_bin_0420 = frame (4k)
frame_vm_group_bin_0421 = frame (4k)
frame_vm_group_bin_0422 = frame (4k)
frame_vm_group_bin_0423 = frame (4k)
frame_vm_group_bin_0424 = frame (4k)
frame_vm_group_bin_0425 = frame (4k)
frame_vm_group_bin_0426 = frame (4k)
frame_vm_group_bin_0427 = frame (4k)
frame_vm_group_bin_0428 = frame (4k)
frame_vm_group_bin_0429 = frame (4k)
frame_vm_group_bin_0430 = frame (4k)
frame_vm_group_bin_0431 = frame (4k)
frame_vm_group_bin_0432 = frame (4k)
frame_vm_group_bin_0433 = frame (4k)
frame_vm_group_bin_0434 = frame (4k)
frame_vm_group_bin_0435 = frame (4k)
frame_vm_group_bin_0436 = frame (4k)
frame_vm_group_bin_0437 = frame (4k)
frame_vm_group_bin_0438 = frame (4k)
frame_vm_group_bin_0439 = frame (4k)
frame_vm_group_bin_0440 = frame (4k)
frame_vm_group_bin_0441 = frame (4k)
frame_vm_group_bin_0442 = frame (4k)
frame_vm_group_bin_0443 = frame (4k)
frame_vm_group_bin_0444 = frame (4k)
frame_vm_group_bin_0445 = frame (4k)
frame_vm_group_bin_0446 = frame (4k)
frame_vm_group_bin_0447 = frame (4k)
frame_vm_group_bin_0448 = frame (4k)
frame_vm_group_bin_0449 = frame (4k)
frame_vm_group_bin_0450 = frame (4k)
frame_vm_group_bin_0451 = frame (4k)
frame_vm_group_bin_0452 = frame (4k)
frame_vm_group_bin_0453 = frame (4k)
frame_vm_group_bin_0454 = frame (4k)
frame_vm_group_bin_0455 = frame (4k)
frame_vm_group_bin_0456 = frame (4k)
frame_vm_group_bin_0457 = frame (4k)
frame_vm_group_bin_0458 = frame (4k)
frame_vm_group_bin_0459 = frame (4k)
frame_vm_group_bin_0460 = frame (4k)
frame_vm_group_bin_0461 = frame (4k)
frame_vm_group_bin_0462 = frame (4k)
frame_vm_group_bin_0463 = frame (4k)
frame_vm_group_bin_0464 = frame (4k)
frame_vm_group_bin_0465 = frame (4k)
frame_vm_group_bin_0466 = frame (4k)
frame_vm_group_bin_0467 = frame (4k)
frame_vm_group_bin_0468 = frame (4k)
frame_vm_group_bin_0469 = frame (4k)
frame_vm_group_bin_0470 = frame (4k)
frame_vm_group_bin_0471 = frame (4k)
frame_vm_group_bin_0472 = frame (4k)
frame_vm_group_bin_0473 = frame (4k)
frame_vm_group_bin_0474 = frame (4k)
frame_vm_group_bin_0475 = frame (4k)
frame_vm_group_bin_0476 = frame (4k)
frame_vm_group_bin_0477 = frame (4k)
frame_vm_group_bin_0478 = frame (4k)
frame_vm_group_bin_0479 = frame (4k)
frame_vm_group_bin_0480 = frame (4k)
frame_vm_group_bin_0481 = frame (4k)
frame_vm_group_bin_0482 = frame (4k)
frame_vm_group_bin_0483 = frame (4k)
frame_vm_group_bin_0484 = frame (4k)
frame_vm_group_bin_0485 = frame (4k)
frame_vm_group_bin_0486 = frame (4k)
frame_vm_group_bin_0487 = frame (4k)
frame_vm_group_bin_0488 = frame (4k)
frame_vm_group_bin_0489 = frame (4k)
frame_vm_group_bin_0490 = frame (4k)
frame_vm_group_bin_0491 = frame (4k)
frame_vm_group_bin_0492 = frame (4k)
frame_vm_group_bin_0493 = frame (4k)
frame_vm_group_bin_0494 = frame (4k)
frame_vm_group_bin_0495 = frame (4k)
frame_vm_group_bin_0496 = frame (4k)
frame_vm_group_bin_0497 = frame (4k)
frame_vm_group_bin_0498 = frame (4k)
frame_vm_group_bin_0499 = frame (4k)
frame_vm_group_bin_0500 = frame (4k)
frame_vm_group_bin_0501 = frame (4k)
frame_vm_group_bin_0502 = frame (4k)
frame_vm_group_bin_0503 = frame (4k)
frame_vm_group_bin_0504 = frame (4k)
frame_vm_group_bin_0505 = frame (4k)
frame_vm_group_bin_0506 = frame (4k)
frame_vm_group_bin_0507 = frame (4k)
frame_vm_group_bin_0508 = frame (4k)
frame_vm_group_bin_0509 = frame (4k)
frame_vm_group_bin_0510 = frame (4k)
frame_vm_group_bin_0511 = frame (4k)
frame_vm_group_bin_0512 = frame (4k)
frame_vm_group_bin_0513 = frame (4k)
frame_vm_group_bin_0514 = frame (4k)
frame_vm_group_bin_0515 = frame (4k)
frame_vm_group_bin_0516 = frame (4k)
frame_vm_group_bin_0517 = frame (4k)
frame_vm_group_bin_0518 = frame (4k)
frame_vm_group_bin_0519 = frame (4k)
frame_vm_group_bin_0520 = frame (4k)
frame_vm_group_bin_0521 = frame (4k)
frame_vm_group_bin_0522 = frame (4k)
frame_vm_group_bin_0523 = frame (4k)
frame_vm_group_bin_0524 = frame (4k)
frame_vm_group_bin_0525 = frame (4k)
frame_vm_group_bin_0526 = frame (4k)
frame_vm_group_bin_0527 = frame (4k)
frame_vm_group_bin_0528 = frame (4k)
frame_vm_group_bin_0529 = frame (4k)
frame_vm_group_bin_0530 = frame (4k)
frame_vm_group_bin_0531 = frame (4k)
frame_vm_group_bin_0532 = frame (4k)
frame_vm_group_bin_0533 = frame (4k)
frame_vm_group_bin_0534 = frame (4k)
frame_vm_group_bin_0535 = frame (4k)
frame_vm_group_bin_0536 = frame (4k)
frame_vm_group_bin_0537 = frame (4k)
frame_vm_group_bin_0538 = frame (4k)
frame_vm_group_bin_0539 = frame (4k)
frame_vm_group_bin_0540 = frame (4k)
frame_vm_group_bin_0541 = frame (4k)
frame_vm_group_bin_0542 = frame (4k)
frame_vm_group_bin_0543 = frame (4k)
frame_vm_group_bin_0544 = frame (4k)
frame_vm_group_bin_0545 = frame (4k)
frame_vm_group_bin_0546 = frame (4k)
frame_vm_group_bin_0547 = frame (4k)
frame_vm_group_bin_0548 = frame (4k)
frame_vm_group_bin_0549 = frame (4k)
frame_vm_group_bin_0550 = frame (4k)
frame_vm_group_bin_0551 = frame (4k)
frame_vm_group_bin_0552 = frame (4k)
frame_vm_group_bin_0553 = frame (4k)
frame_vm_group_bin_0554 = frame (4k)
frame_vm_group_bin_0555 = frame (4k)
frame_vm_group_bin_0556 = frame (4k)
frame_vm_group_bin_0557 = frame (4k)
frame_vm_group_bin_0558 = frame (4k)
frame_vm_group_bin_0559 = frame (4k)
frame_vm_group_bin_0560 = frame (4k)
frame_vm_group_bin_0561 = frame (4k)
frame_vm_group_bin_0562 = frame (4k)
frame_vm_group_bin_0563 = frame (4k)
frame_vm_group_bin_0564 = frame (4k)
frame_vm_group_bin_0565 = frame (4k)
frame_vm_group_bin_0566 = frame (4k)
frame_vm_group_bin_0567 = frame (4k)
frame_vm_group_bin_0568 = frame (4k)
frame_vm_group_bin_0569 = frame (4k)
frame_vm_group_bin_0570 = frame (4k)
frame_vm_group_bin_0571 = frame (4k)
frame_vm_group_bin_0572 = frame (4k)
frame_vm_group_bin_0573 = frame (4k)
frame_vm_group_bin_0574 = frame (4k)
frame_vm_group_bin_0575 = frame (4k)
frame_vm_group_bin_0576 = frame (4k)
frame_vm_group_bin_0577 = frame (4k)
frame_vm_group_bin_0578 = frame (4k)
frame_vm_group_bin_0579 = frame (4k)
frame_vm_group_bin_0580 = frame (4k)
frame_vm_group_bin_0581 = frame (4k)
frame_vm_group_bin_0582 = frame (4k)
frame_vm_group_bin_0583 = frame (4k)
frame_vm_group_bin_0584 = frame (4k)
frame_vm_group_bin_0585 = frame (4k)
frame_vm_group_bin_0586 = frame (4k)
frame_vm_group_bin_0587 = frame (4k)
frame_vm_group_bin_0588 = frame (4k)
frame_vm_group_bin_0589 = frame (4k)
frame_vm_group_bin_0590 = frame (4k)
frame_vm_group_bin_0591 = frame (4k)
frame_vm_group_bin_0592 = frame (4k)
frame_vm_group_bin_0593 = frame (4k)
frame_vm_group_bin_0594 = frame (4k)
frame_vm_group_bin_0595 = frame (4k)
frame_vm_group_bin_0596 = frame (4k)
frame_vm_group_bin_0597 = frame (4k)
frame_vm_group_bin_0598 = frame (4k)
frame_vm_group_bin_0599 = frame (4k)
frame_vm_group_bin_0600 = frame (4k)
frame_vm_group_bin_0601 = frame (4k)
frame_vm_group_bin_0602 = frame (4k)
frame_vm_group_bin_0603 = frame (4k)
frame_vm_group_bin_0604 = frame (4k)
frame_vm_group_bin_0605 = frame (4k)
frame_vm_group_bin_0606 = frame (4k)
frame_vm_group_bin_0607 = frame (4k)
frame_vm_group_bin_0608 = frame (4k)
frame_vm_group_bin_0609 = frame (4k)
frame_vm_group_bin_0610 = frame (4k)
frame_vm_group_bin_0611 = frame (4k)
frame_vm_group_bin_0612 = frame (4k)
frame_vm_group_bin_0613 = frame (4k)
frame_vm_group_bin_0614 = frame (4k)
frame_vm_group_bin_0615 = frame (4k)
frame_vm_group_bin_0616 = frame (4k)
frame_vm_group_bin_0617 = frame (4k)
frame_vm_group_bin_0618 = frame (4k)
frame_vm_group_bin_0619 = frame (4k)
frame_vm_group_bin_0620 = frame (4k)
frame_vm_group_bin_0621 = frame (4k)
frame_vm_group_bin_0622 = frame (4k)
frame_vm_group_bin_0623 = frame (4k)
frame_vm_group_bin_0624 = frame (4k)
frame_vm_group_bin_0625 = frame (4k)
frame_vm_group_bin_0626 = frame (4k)
frame_vm_group_bin_0627 = frame (4k)
frame_vm_group_bin_0628 = frame (4k)
frame_vm_group_bin_0629 = frame (4k)
frame_vm_group_bin_0630 = frame (4k)
frame_vm_group_bin_0631 = frame (4k)
frame_vm_group_bin_0632 = frame (4k)
frame_vm_group_bin_0633 = frame (4k)
frame_vm_group_bin_0634 = frame (4k)
frame_vm_group_bin_0635 = frame (4k)
frame_vm_group_bin_0636 = frame (4k)
frame_vm_group_bin_0637 = frame (4k)
frame_vm_group_bin_0638 = frame (4k)
frame_vm_group_bin_0639 = frame (4k)
frame_vm_group_bin_0640 = frame (4k)
frame_vm_group_bin_0641 = frame (4k)
frame_vm_group_bin_0642 = frame (4k)
frame_vm_group_bin_0643 = frame (4k)
frame_vm_group_bin_0644 = frame (4k)
frame_vm_group_bin_0645 = frame (4k)
frame_vm_group_bin_0646 = frame (4k)
frame_vm_group_bin_0647 = frame (4k)
frame_vm_group_bin_0648 = frame (4k)
frame_vm_group_bin_0649 = frame (4k)
frame_vm_group_bin_0650 = frame (4k)
frame_vm_group_bin_0651 = frame (4k)
frame_vm_group_bin_0652 = frame (4k)
frame_vm_group_bin_0653 = frame (4k)
frame_vm_group_bin_0654 = frame (4k)
frame_vm_group_bin_0655 = frame (4k)
frame_vm_group_bin_0656 = frame (4k)
frame_vm_group_bin_0657 = frame (4k)
frame_vm_group_bin_0658 = frame (4k)
frame_vm_group_bin_0659 = frame (4k)
frame_vm_group_bin_0660 = frame (4k)
frame_vm_group_bin_0661 = frame (4k)
frame_vm_group_bin_0662 = frame (4k)
frame_vm_group_bin_0663 = frame (4k)
frame_vm_group_bin_0664 = frame (4k)
frame_vm_group_bin_0665 = frame (4k)
frame_vm_group_bin_0666 = frame (4k)
frame_vm_group_bin_0667 = frame (4k)
frame_vm_group_bin_0668 = frame (4k)
frame_vm_group_bin_0669 = frame (4k)
frame_vm_group_bin_0670 = frame (4k)
frame_vm_group_bin_0671 = frame (4k)
frame_vm_group_bin_0672 = frame (4k)
frame_vm_group_bin_0673 = frame (4k)
frame_vm_group_bin_0674 = frame (4k)
frame_vm_group_bin_0675 = frame (4k)
frame_vm_group_bin_0676 = frame (4k)
frame_vm_group_bin_0677 = frame (4k)
frame_vm_group_bin_0678 = frame (4k)
frame_vm_group_bin_0679 = frame (4k)
frame_vm_group_bin_0680 = frame (4k)
frame_vm_group_bin_0681 = frame (4k)
frame_vm_group_bin_0682 = frame (4k)
frame_vm_group_bin_0683 = frame (4k)
frame_vm_group_bin_0684 = frame (4k)
frame_vm_group_bin_0685 = frame (4k)
frame_vm_group_bin_0686 = frame (4k)
frame_vm_group_bin_0687 = frame (4k)
frame_vm_group_bin_0688 = frame (4k)
frame_vm_group_bin_0689 = frame (4k)
frame_vm_group_bin_0690 = frame (4k)
frame_vm_group_bin_0691 = frame (4k)
frame_vm_group_bin_0692 = frame (4k)
frame_vm_group_bin_0693 = frame (4k)
frame_vm_group_bin_0694 = frame (4k)
frame_vm_group_bin_0695 = frame (4k)
frame_vm_group_bin_0696 = frame (4k)
frame_vm_group_bin_0697 = frame (4k)
frame_vm_group_bin_0698 = frame (4k)
frame_vm_group_bin_0699 = frame (4k)
frame_vm_group_bin_0700 = frame (4k)
frame_vm_group_bin_0701 = frame (4k)
frame_vm_group_bin_0702 = frame (4k)
frame_vm_group_bin_0703 = frame (4k)
frame_vm_group_bin_0704 = frame (4k)
frame_vm_group_bin_0705 = frame (4k)
frame_vm_group_bin_0706 = frame (4k)
frame_vm_group_bin_0707 = frame (4k)
frame_vm_group_bin_0708 = frame (4k)
frame_vm_group_bin_0709 = frame (4k)
frame_vm_group_bin_0710 = frame (4k)
frame_vm_group_bin_0711 = frame (4k)
frame_vm_group_bin_0712 = frame (4k)
frame_vm_group_bin_0713 = frame (4k)
frame_vm_group_bin_0714 = frame (4k)
frame_vm_group_bin_0715 = frame (4k)
frame_vm_group_bin_0716 = frame (4k)
frame_vm_group_bin_0717 = frame (4k)
frame_vm_group_bin_0718 = frame (4k)
frame_vm_group_bin_0719 = frame (4k)
frame_vm_group_bin_0720 = frame (4k)
frame_vm_group_bin_0721 = frame (4k)
frame_vm_group_bin_0722 = frame (4k)
frame_vm_group_bin_0723 = frame (4k)
frame_vm_group_bin_0724 = frame (4k)
frame_vm_group_bin_0725 = frame (4k)
frame_vm_group_bin_0726 = frame (4k)
frame_vm_group_bin_0727 = frame (4k)
frame_vm_group_bin_0728 = frame (4k)
frame_vm_group_bin_0729 = frame (4k)
frame_vm_group_bin_0730 = frame (4k)
frame_vm_group_bin_0731 = frame (4k)
frame_vm_group_bin_0732 = frame (4k)
frame_vm_group_bin_0733 = frame (4k)
frame_vm_group_bin_0734 = frame (4k)
frame_vm_group_bin_0735 = frame (4k)
frame_vm_group_bin_0736 = frame (4k)
frame_vm_group_bin_0737 = frame (4k)
frame_vm_group_bin_0738 = frame (4k)
frame_vm_group_bin_0739 = frame (4k)
frame_vm_group_bin_0740 = frame (4k)
frame_vm_group_bin_0741 = frame (4k)
frame_vm_group_bin_0742 = frame (4k)
frame_vm_group_bin_0743 = frame (4k)
frame_vm_group_bin_0744 = frame (4k)
frame_vm_group_bin_0745 = frame (4k)
frame_vm_group_bin_0746 = frame (4k)
frame_vm_group_bin_0747 = frame (4k)
frame_vm_group_bin_0748 = frame (4k)
frame_vm_group_bin_0749 = frame (4k)
frame_vm_group_bin_0750 = frame (4k)
frame_vm_group_bin_0751 = frame (4k)
frame_vm_group_bin_0752 = frame (4k)
frame_vm_group_bin_0753 = frame (4k)
frame_vm_group_bin_0754 = frame (4k)
frame_vm_group_bin_0755 = frame (4k)
frame_vm_group_bin_0756 = frame (4k)
frame_vm_group_bin_0757 = frame (4k)
frame_vm_group_bin_0758 = frame (4k)
frame_vm_group_bin_0759 = frame (4k)
frame_vm_group_bin_0760 = frame (4k)
frame_vm_group_bin_0761 = frame (4k)
frame_vm_group_bin_0762 = frame (4k)
frame_vm_group_bin_0763 = frame (4k)
frame_vm_group_bin_0764 = frame (4k)
frame_vm_group_bin_0765 = frame (4k)
frame_vm_group_bin_0766 = frame (4k)
frame_vm_group_bin_0767 = frame (4k)
frame_vm_group_bin_0768 = frame (4k)
frame_vm_group_bin_0769 = frame (4k)
frame_vm_group_bin_0770 = frame (4k)
frame_vm_group_bin_0771 = frame (4k)
frame_vm_group_bin_0772 = frame (4k)
frame_vm_group_bin_0773 = frame (4k)
frame_vm_group_bin_0774 = frame (4k)
frame_vm_group_bin_0775 = frame (4k)
frame_vm_group_bin_0776 = frame (4k)
frame_vm_group_bin_0777 = frame (4k)
frame_vm_group_bin_0778 = frame (4k)
frame_vm_group_bin_0779 = frame (4k)
frame_vm_group_bin_0780 = frame (4k)
frame_vm_group_bin_0781 = frame (4k)
frame_vm_group_bin_0782 = frame (4k)
frame_vm_group_bin_0783 = frame (4k)
frame_vm_group_bin_0784 = frame (4k)
frame_vm_group_bin_0785 = frame (4k)
frame_vm_group_bin_0786 = frame (4k)
frame_vm_group_bin_0787 = frame (4k)
frame_vm_group_bin_0788 = frame (4k)
frame_vm_group_bin_0789 = frame (4k)
frame_vm_group_bin_0790 = frame (4k)
frame_vm_group_bin_0791 = frame (4k)
frame_vm_group_bin_0792 = frame (4k)
frame_vm_group_bin_0793 = frame (4k)
frame_vm_group_bin_0794 = frame (4k)
frame_vm_group_bin_0795 = frame (4k)
frame_vm_group_bin_0796 = frame (4k)
frame_vm_group_bin_0797 = frame (4k)
frame_vm_group_bin_0798 = frame (4k)
frame_vm_group_bin_0799 = frame (4k)
frame_vm_group_bin_0800 = frame (4k)
frame_vm_group_bin_0801 = frame (4k)
frame_vm_group_bin_0802 = frame (4k)
frame_vm_group_bin_0803 = frame (4k)
frame_vm_group_bin_0804 = frame (4k)
frame_vm_group_bin_0805 = frame (4k)
frame_vm_group_bin_0806 = frame (4k)
frame_vm_group_bin_0807 = frame (4k)
frame_vm_group_bin_0808 = frame (4k)
frame_vm_group_bin_0809 = frame (4k)
frame_vm_group_bin_0810 = frame (4k)
frame_vm_group_bin_0811 = frame (4k)
frame_vm_group_bin_0812 = frame (4k)
frame_vm_group_bin_0813 = frame (4k)
frame_vm_group_bin_0814 = frame (4k)
frame_vm_group_bin_0815 = frame (4k)
frame_vm_group_bin_0816 = frame (4k)
frame_vm_group_bin_0817 = frame (4k)
frame_vm_group_bin_0818 = frame (4k)
frame_vm_group_bin_0819 = frame (4k)
frame_vm_group_bin_0820 = frame (4k)
frame_vm_group_bin_0821 = frame (4k)
frame_vm_group_bin_0822 = frame (4k)
frame_vm_group_bin_0823 = frame (4k)
frame_vm_group_bin_0824 = frame (4k)
frame_vm_group_bin_0825 = frame (4k)
frame_vm_group_bin_0826 = frame (4k)
frame_vm_group_bin_0827 = frame (4k)
frame_vm_group_bin_0828 = frame (4k)
frame_vm_group_bin_0829 = frame (4k)
frame_vm_group_bin_0830 = frame (4k)
frame_vm_group_bin_0831 = frame (4k)
frame_vm_group_bin_0832 = frame (4k)
frame_vm_group_bin_0833 = frame (4k)
frame_vm_group_bin_0834 = frame (4k)
frame_vm_group_bin_0835 = frame (4k)
frame_vm_group_bin_0836 = frame (4k)
frame_vm_group_bin_0837 = frame (4k)
frame_vm_group_bin_0838 = frame (4k)
frame_vm_group_bin_0839 = frame (4k)
frame_vm_group_bin_0840 = frame (4k)
frame_vm_group_bin_0841 = frame (4k)
frame_vm_group_bin_0842 = frame (4k)
frame_vm_group_bin_0843 = frame (4k)
frame_vm_group_bin_0844 = frame (4k)
frame_vm_group_bin_0845 = frame (4k)
frame_vm_group_bin_0846 = frame (4k)
frame_vm_group_bin_0847 = frame (4k)
frame_vm_group_bin_0848 = frame (4k)
frame_vm_group_bin_0849 = frame (4k)
frame_vm_group_bin_0850 = frame (4k)
frame_vm_group_bin_0851 = frame (4k)
frame_vm_group_bin_0852 = frame (4k)
frame_vm_group_bin_0853 = frame (4k)
frame_vm_group_bin_0854 = frame (4k)
frame_vm_group_bin_0855 = frame (4k)
frame_vm_group_bin_0856 = frame (4k)
frame_vm_group_bin_0857 = frame (4k)
frame_vm_group_bin_0858 = frame (4k)
frame_vm_group_bin_0859 = frame (4k)
frame_vm_group_bin_0860 = frame (4k)
frame_vm_group_bin_0861 = frame (4k)
frame_vm_group_bin_0862 = frame (4k)
frame_vm_group_bin_0863 = frame (4k)
frame_vm_group_bin_0864 = frame (4k)
frame_vm_group_bin_0865 = frame (4k)
frame_vm_group_bin_0866 = frame (4k)
frame_vm_group_bin_0867 = frame (4k)
frame_vm_group_bin_0868 = frame (4k)
frame_vm_group_bin_0869 = frame (4k)
frame_vm_group_bin_0870 = frame (4k)
frame_vm_group_bin_0871 = frame (4k)
frame_vm_group_bin_0872 = frame (4k)
frame_vm_group_bin_0873 = frame (4k)
frame_vm_group_bin_0874 = frame (4k)
frame_vm_group_bin_0875 = frame (4k)
frame_vm_group_bin_0876 = frame (4k)
frame_vm_group_bin_0877 = frame (4k)
frame_vm_group_bin_0878 = frame (4k)
frame_vm_group_bin_0879 = frame (4k)
frame_vm_group_bin_0880 = frame (4k)
frame_vm_group_bin_0881 = frame (4k)
frame_vm_group_bin_0882 = frame (4k)
frame_vm_group_bin_0883 = frame (4k)
frame_vm_group_bin_0884 = frame (4k)
frame_vm_group_bin_0885 = frame (4k)
frame_vm_group_bin_0886 = frame (4k)
frame_vm_group_bin_0887 = frame (4k)
frame_vm_group_bin_0888 = frame (4k)
frame_vm_group_bin_0889 = frame (4k)
frame_vm_group_bin_0890 = frame (4k)
frame_vm_group_bin_0891 = frame (4k)
frame_vm_group_bin_0892 = frame (4k)
frame_vm_group_bin_0893 = frame (4k)
frame_vm_group_bin_0894 = frame (4k)
frame_vm_group_bin_0895 = frame (4k)
frame_vm_group_bin_0896 = frame (4k)
frame_vm_group_bin_0897 = frame (4k)
frame_vm_group_bin_0898 = frame (4k)
frame_vm_group_bin_0899 = frame (4k)
frame_vm_group_bin_0900 = frame (4k)
frame_vm_group_bin_0901 = frame (4k)
frame_vm_group_bin_0902 = frame (4k)
frame_vm_group_bin_0903 = frame (4k)
frame_vm_group_bin_0904 = frame (4k)
frame_vm_group_bin_0905 = frame (4k)
frame_vm_group_bin_0906 = frame (4k)
frame_vm_group_bin_0907 = frame (4k)
frame_vm_group_bin_0908 = frame (4k)
frame_vm_group_bin_0909 = frame (4k)
frame_vm_group_bin_0910 = frame (4k)
frame_vm_group_bin_0911 = frame (4k)
frame_vm_group_bin_0912 = frame (4k)
frame_vm_group_bin_0913 = frame (4k)
frame_vm_group_bin_0914 = frame (4k)
frame_vm_group_bin_0915 = frame (4k)
frame_vm_group_bin_0916 = frame (4k)
frame_vm_group_bin_0917 = frame (4k)
frame_vm_group_bin_0918 = frame (4k)
frame_vm_group_bin_0919 = frame (4k)
frame_vm_group_bin_0920 = frame (4k)
frame_vm_group_bin_0921 = frame (4k)
frame_vm_group_bin_0922 = frame (4k)
frame_vm_group_bin_0923 = frame (4k)
frame_vm_group_bin_0924 = frame (4k)
frame_vm_group_bin_0925 = frame (4k)
frame_vm_group_bin_0926 = frame (4k)
frame_vm_group_bin_0927 = frame (4k)
frame_vm_group_bin_0928 = frame (4k)
frame_vm_group_bin_0929 = frame (4k)
frame_vm_group_bin_0930 = frame (4k)
frame_vm_group_bin_0931 = frame (4k)
frame_vm_group_bin_0932 = frame (4k)
frame_vm_group_bin_0933 = frame (4k)
frame_vm_group_bin_0934 = frame (4k)
frame_vm_group_bin_0935 = frame (4k)
frame_vm_group_bin_0936 = frame (4k)
frame_vm_group_bin_0937 = frame (4k)
frame_vm_group_bin_0938 = frame (4k)
frame_vm_group_bin_0939 = frame (4k)
frame_vm_group_bin_0940 = frame (4k)
frame_vm_group_bin_0941 = frame (4k)
frame_vm_group_bin_0942 = frame (4k)
frame_vm_group_bin_0943 = frame (4k)
frame_vm_group_bin_0944 = frame (4k)
frame_vm_group_bin_0945 = frame (4k)
frame_vm_group_bin_0946 = frame (4k)
frame_vm_group_bin_0947 = frame (4k)
frame_vm_group_bin_0948 = frame (4k)
frame_vm_group_bin_0949 = frame (4k)
frame_vm_group_bin_0950 = frame (4k)
frame_vm_group_bin_0951 = frame (4k)
frame_vm_group_bin_0952 = frame (4k)
frame_vm_group_bin_0953 = frame (4k)
frame_vm_group_bin_0954 = frame (4k)
frame_vm_group_bin_0955 = frame (4k)
frame_vm_group_bin_0956 = frame (4k)
frame_vm_group_bin_0957 = frame (4k)
frame_vm_group_bin_0958 = frame (4k)
frame_vm_group_bin_0959 = frame (4k)
frame_vm_group_bin_0960 = frame (4k)
frame_vm_group_bin_0961 = frame (4k)
frame_vm_group_bin_0962 = frame (4k)
frame_vm_group_bin_0963 = frame (4k)
frame_vm_group_bin_0964 = frame (4k)
frame_vm_group_bin_0965 = frame (4k)
frame_vm_group_bin_0966 = frame (4k)
frame_vm_group_bin_0967 = frame (4k)
frame_vm_group_bin_0968 = frame (4k)
frame_vm_group_bin_0969 = frame (4k)
frame_vm_group_bin_0970 = frame (4k)
frame_vm_group_bin_0971 = frame (4k)
frame_vm_group_bin_0972 = frame (4k)
frame_vm_group_bin_0973 = frame (4k)
frame_vm_group_bin_0974 = frame (4k)
frame_vm_group_bin_0975 = frame (4k)
frame_vm_group_bin_0976 = frame (4k)
frame_vm_group_bin_0977 = frame (4k)
frame_vm_group_bin_0978 = frame (4k)
frame_vm_group_bin_0979 = frame (4k)
frame_vm_group_bin_0980 = frame (4k)
frame_vm_group_bin_0981 = frame (4k)
frame_vm_group_bin_0982 = frame (4k)
frame_vm_group_bin_0983 = frame (4k)
frame_vm_group_bin_0984 = frame (4k)
frame_vm_group_bin_0985 = frame (4k)
frame_vm_group_bin_0986 = frame (4k)
frame_vm_group_bin_0987 = frame (4k)
frame_vm_group_bin_0988 = frame (4k)
frame_vm_group_bin_0989 = frame (4k)
frame_vm_group_bin_0990 = frame (4k)
frame_vm_group_bin_0991 = frame (4k)
frame_vm_group_bin_0992 = frame (4k)
frame_vm_group_bin_0993 = frame (4k)
frame_vm_group_bin_0994 = frame (4k)
frame_vm_group_bin_0995 = frame (4k)
frame_vm_group_bin_0996 = frame (4k)
frame_vm_group_bin_0997 = frame (4k)
frame_vm_group_bin_0998 = frame (4k)
frame_vm_group_bin_0999 = frame (4k)
frame_vm_group_bin_1000 = frame (4k)
frame_vm_group_bin_10000 = frame (4k)
frame_vm_group_bin_10001 = frame (4k)
frame_vm_group_bin_10002 = frame (4k)
frame_vm_group_bin_10003 = frame (4k)
frame_vm_group_bin_10004 = frame (4k)
frame_vm_group_bin_10005 = frame (4k)
frame_vm_group_bin_10006 = frame (4k)
frame_vm_group_bin_10007 = frame (4k)
frame_vm_group_bin_10008 = frame (4k)
frame_vm_group_bin_10009 = frame (4k)
frame_vm_group_bin_1001 = frame (4k)
frame_vm_group_bin_10010 = frame (4k)
frame_vm_group_bin_10011 = frame (4k)
frame_vm_group_bin_10012 = frame (4k)
frame_vm_group_bin_10013 = frame (4k)
frame_vm_group_bin_10014 = frame (4k)
frame_vm_group_bin_10015 = frame (4k)
frame_vm_group_bin_10016 = frame (4k)
frame_vm_group_bin_10017 = frame (4k)
frame_vm_group_bin_10018 = frame (4k)
frame_vm_group_bin_10019 = frame (4k)
frame_vm_group_bin_1002 = frame (4k)
frame_vm_group_bin_10020 = frame (4k)
frame_vm_group_bin_10021 = frame (4k)
frame_vm_group_bin_10022 = frame (4k)
frame_vm_group_bin_10023 = frame (4k)
frame_vm_group_bin_10024 = frame (4k)
frame_vm_group_bin_10025 = frame (4k)
frame_vm_group_bin_10026 = frame (4k)
frame_vm_group_bin_10027 = frame (4k)
frame_vm_group_bin_10028 = frame (4k)
frame_vm_group_bin_10029 = frame (4k)
frame_vm_group_bin_1003 = frame (4k)
frame_vm_group_bin_10030 = frame (4k)
frame_vm_group_bin_10031 = frame (4k)
frame_vm_group_bin_10032 = frame (4k)
frame_vm_group_bin_10033 = frame (4k)
frame_vm_group_bin_10034 = frame (4k)
frame_vm_group_bin_10035 = frame (4k)
frame_vm_group_bin_10036 = frame (4k)
frame_vm_group_bin_10037 = frame (4k)
frame_vm_group_bin_10038 = frame (4k)
frame_vm_group_bin_10039 = frame (4k)
frame_vm_group_bin_1004 = frame (4k)
frame_vm_group_bin_10040 = frame (4k)
frame_vm_group_bin_10041 = frame (4k)
frame_vm_group_bin_10042 = frame (4k)
frame_vm_group_bin_10043 = frame (4k)
frame_vm_group_bin_10044 = frame (4k)
frame_vm_group_bin_10045 = frame (4k)
frame_vm_group_bin_10046 = frame (4k)
frame_vm_group_bin_10047 = frame (4k)
frame_vm_group_bin_10048 = frame (4k)
frame_vm_group_bin_10049 = frame (4k)
frame_vm_group_bin_1005 = frame (4k)
frame_vm_group_bin_10050 = frame (4k)
frame_vm_group_bin_10051 = frame (4k)
frame_vm_group_bin_10052 = frame (4k)
frame_vm_group_bin_10053 = frame (4k)
frame_vm_group_bin_10054 = frame (4k)
frame_vm_group_bin_10055 = frame (4k)
frame_vm_group_bin_10056 = frame (4k)
frame_vm_group_bin_10057 = frame (4k)
frame_vm_group_bin_10058 = frame (4k)
frame_vm_group_bin_10059 = frame (4k)
frame_vm_group_bin_1006 = frame (4k)
frame_vm_group_bin_10060 = frame (4k)
frame_vm_group_bin_10061 = frame (4k)
frame_vm_group_bin_10062 = frame (4k)
frame_vm_group_bin_10063 = frame (4k)
frame_vm_group_bin_10064 = frame (4k)
frame_vm_group_bin_10065 = frame (4k)
frame_vm_group_bin_10066 = frame (4k)
frame_vm_group_bin_10067 = frame (4k)
frame_vm_group_bin_10068 = frame (4k)
frame_vm_group_bin_10069 = frame (4k)
frame_vm_group_bin_1007 = frame (4k)
frame_vm_group_bin_10070 = frame (4k)
frame_vm_group_bin_10071 = frame (4k)
frame_vm_group_bin_10072 = frame (4k)
frame_vm_group_bin_10073 = frame (4k)
frame_vm_group_bin_10074 = frame (4k)
frame_vm_group_bin_10075 = frame (4k)
frame_vm_group_bin_10076 = frame (4k)
frame_vm_group_bin_10077 = frame (4k)
frame_vm_group_bin_10078 = frame (4k)
frame_vm_group_bin_10079 = frame (4k)
frame_vm_group_bin_1008 = frame (4k)
frame_vm_group_bin_10080 = frame (4k)
frame_vm_group_bin_10081 = frame (4k)
frame_vm_group_bin_10082 = frame (4k)
frame_vm_group_bin_10083 = frame (4k)
frame_vm_group_bin_10084 = frame (4k)
frame_vm_group_bin_10085 = frame (4k)
frame_vm_group_bin_10086 = frame (4k)
frame_vm_group_bin_10087 = frame (4k)
frame_vm_group_bin_10088 = frame (4k)
frame_vm_group_bin_10089 = frame (4k)
frame_vm_group_bin_1009 = frame (4k)
frame_vm_group_bin_10090 = frame (4k)
frame_vm_group_bin_10091 = frame (4k)
frame_vm_group_bin_10092 = frame (4k)
frame_vm_group_bin_10093 = frame (4k)
frame_vm_group_bin_10094 = frame (4k)
frame_vm_group_bin_10095 = frame (4k)
frame_vm_group_bin_10096 = frame (4k)
frame_vm_group_bin_10097 = frame (4k)
frame_vm_group_bin_10098 = frame (4k)
frame_vm_group_bin_10099 = frame (4k)
frame_vm_group_bin_1010 = frame (4k)
frame_vm_group_bin_10100 = frame (4k)
frame_vm_group_bin_10101 = frame (4k)
frame_vm_group_bin_10102 = frame (4k)
frame_vm_group_bin_10103 = frame (4k)
frame_vm_group_bin_10104 = frame (4k)
frame_vm_group_bin_10105 = frame (4k)
frame_vm_group_bin_10106 = frame (4k)
frame_vm_group_bin_10107 = frame (4k)
frame_vm_group_bin_10108 = frame (4k)
frame_vm_group_bin_10109 = frame (4k)
frame_vm_group_bin_1011 = frame (4k)
frame_vm_group_bin_10110 = frame (4k)
frame_vm_group_bin_10111 = frame (4k)
frame_vm_group_bin_10112 = frame (4k)
frame_vm_group_bin_10113 = frame (4k)
frame_vm_group_bin_10114 = frame (4k)
frame_vm_group_bin_10115 = frame (4k)
frame_vm_group_bin_10116 = frame (4k)
frame_vm_group_bin_10117 = frame (4k)
frame_vm_group_bin_10118 = frame (4k)
frame_vm_group_bin_10119 = frame (4k)
frame_vm_group_bin_1012 = frame (4k)
frame_vm_group_bin_10120 = frame (4k)
frame_vm_group_bin_10121 = frame (4k)
frame_vm_group_bin_10122 = frame (4k)
frame_vm_group_bin_10123 = frame (4k)
frame_vm_group_bin_10124 = frame (4k)
frame_vm_group_bin_10125 = frame (4k)
frame_vm_group_bin_10126 = frame (4k)
frame_vm_group_bin_10127 = frame (4k)
frame_vm_group_bin_10128 = frame (4k)
frame_vm_group_bin_10129 = frame (4k)
frame_vm_group_bin_1013 = frame (4k)
frame_vm_group_bin_10130 = frame (4k)
frame_vm_group_bin_10131 = frame (4k)
frame_vm_group_bin_10132 = frame (4k)
frame_vm_group_bin_10133 = frame (4k)
frame_vm_group_bin_10134 = frame (4k)
frame_vm_group_bin_10135 = frame (4k)
frame_vm_group_bin_10136 = frame (4k)
frame_vm_group_bin_10137 = frame (4k)
frame_vm_group_bin_10138 = frame (4k)
frame_vm_group_bin_10139 = frame (4k)
frame_vm_group_bin_1014 = frame (4k)
frame_vm_group_bin_10140 = frame (4k)
frame_vm_group_bin_10141 = frame (4k)
frame_vm_group_bin_10142 = frame (4k)
frame_vm_group_bin_10143 = frame (4k)
frame_vm_group_bin_10144 = frame (4k)
frame_vm_group_bin_10145 = frame (4k)
frame_vm_group_bin_10146 = frame (4k)
frame_vm_group_bin_10147 = frame (4k)
frame_vm_group_bin_10148 = frame (4k)
frame_vm_group_bin_10149 = frame (4k)
frame_vm_group_bin_1015 = frame (4k)
frame_vm_group_bin_10150 = frame (4k)
frame_vm_group_bin_10151 = frame (4k)
frame_vm_group_bin_10152 = frame (4k)
frame_vm_group_bin_10153 = frame (4k)
frame_vm_group_bin_10154 = frame (4k)
frame_vm_group_bin_10155 = frame (4k)
frame_vm_group_bin_10156 = frame (4k)
frame_vm_group_bin_10157 = frame (4k)
frame_vm_group_bin_10158 = frame (4k)
frame_vm_group_bin_10159 = frame (4k)
frame_vm_group_bin_1016 = frame (4k)
frame_vm_group_bin_10160 = frame (4k)
frame_vm_group_bin_10161 = frame (4k)
frame_vm_group_bin_10162 = frame (4k)
frame_vm_group_bin_10163 = frame (4k)
frame_vm_group_bin_10164 = frame (4k)
frame_vm_group_bin_10165 = frame (4k)
frame_vm_group_bin_10166 = frame (4k)
frame_vm_group_bin_10167 = frame (4k)
frame_vm_group_bin_10168 = frame (4k)
frame_vm_group_bin_10169 = frame (4k)
frame_vm_group_bin_1017 = frame (4k)
frame_vm_group_bin_10170 = frame (4k)
frame_vm_group_bin_10171 = frame (4k)
frame_vm_group_bin_10172 = frame (4k)
frame_vm_group_bin_10173 = frame (4k)
frame_vm_group_bin_10174 = frame (4k)
frame_vm_group_bin_10175 = frame (4k)
frame_vm_group_bin_10176 = frame (4k)
frame_vm_group_bin_10177 = frame (4k)
frame_vm_group_bin_10178 = frame (4k)
frame_vm_group_bin_10179 = frame (4k)
frame_vm_group_bin_1018 = frame (4k)
frame_vm_group_bin_10180 = frame (4k)
frame_vm_group_bin_10181 = frame (4k)
frame_vm_group_bin_10182 = frame (4k)
frame_vm_group_bin_10183 = frame (4k)
frame_vm_group_bin_10184 = frame (4k)
frame_vm_group_bin_10185 = frame (4k)
frame_vm_group_bin_10186 = frame (4k)
frame_vm_group_bin_10187 = frame (4k)
frame_vm_group_bin_10188 = frame (4k)
frame_vm_group_bin_10189 = frame (4k)
frame_vm_group_bin_1019 = frame (4k)
frame_vm_group_bin_10190 = frame (4k)
frame_vm_group_bin_10191 = frame (4k)
frame_vm_group_bin_10192 = frame (4k)
frame_vm_group_bin_10193 = frame (4k)
frame_vm_group_bin_10194 = frame (4k)
frame_vm_group_bin_10195 = frame (4k)
frame_vm_group_bin_10196 = frame (4k)
frame_vm_group_bin_10197 = frame (4k)
frame_vm_group_bin_10198 = frame (4k)
frame_vm_group_bin_10199 = frame (4k)
frame_vm_group_bin_1020 = frame (4k)
frame_vm_group_bin_10200 = frame (4k)
frame_vm_group_bin_10201 = frame (4k)
frame_vm_group_bin_10202 = frame (4k)
frame_vm_group_bin_10203 = frame (4k)
frame_vm_group_bin_10204 = frame (4k)
frame_vm_group_bin_10205 = frame (4k)
frame_vm_group_bin_10206 = frame (4k)
frame_vm_group_bin_10207 = frame (4k)
frame_vm_group_bin_10208 = frame (4k)
frame_vm_group_bin_10209 = frame (4k)
frame_vm_group_bin_1021 = frame (4k)
frame_vm_group_bin_10210 = frame (4k)
frame_vm_group_bin_10211 = frame (4k)
frame_vm_group_bin_10212 = frame (4k)
frame_vm_group_bin_10213 = frame (4k)
frame_vm_group_bin_10214 = frame (4k)
frame_vm_group_bin_10215 = frame (4k)
frame_vm_group_bin_10216 = frame (4k)
frame_vm_group_bin_10217 = frame (4k)
frame_vm_group_bin_10218 = frame (4k)
frame_vm_group_bin_10219 = frame (4k)
frame_vm_group_bin_1022 = frame (4k)
frame_vm_group_bin_10220 = frame (4k)
frame_vm_group_bin_10221 = frame (4k)
frame_vm_group_bin_10222 = frame (4k)
frame_vm_group_bin_10223 = frame (4k)
frame_vm_group_bin_10224 = frame (4k)
frame_vm_group_bin_10225 = frame (4k)
frame_vm_group_bin_10226 = frame (4k)
frame_vm_group_bin_10227 = frame (4k)
frame_vm_group_bin_10228 = frame (4k)
frame_vm_group_bin_10229 = frame (4k)
frame_vm_group_bin_1023 = frame (4k)
frame_vm_group_bin_10230 = frame (4k)
frame_vm_group_bin_10231 = frame (4k)
frame_vm_group_bin_10232 = frame (4k)
frame_vm_group_bin_10233 = frame (4k)
frame_vm_group_bin_10234 = frame (4k)
frame_vm_group_bin_10235 = frame (4k)
frame_vm_group_bin_10236 = frame (4k)
frame_vm_group_bin_10237 = frame (4k)
frame_vm_group_bin_10238 = frame (4k)
frame_vm_group_bin_10239 = frame (4k)
frame_vm_group_bin_1024 = frame (4k)
frame_vm_group_bin_10240 = frame (4k)
frame_vm_group_bin_10241 = frame (4k)
frame_vm_group_bin_10242 = frame (4k)
frame_vm_group_bin_10243 = frame (4k)
frame_vm_group_bin_10244 = frame (4k)
frame_vm_group_bin_10245 = frame (4k)
frame_vm_group_bin_10246 = frame (4k)
frame_vm_group_bin_10247 = frame (4k)
frame_vm_group_bin_10248 = frame (4k)
frame_vm_group_bin_10249 = frame (4k)
frame_vm_group_bin_1025 = frame (4k)
frame_vm_group_bin_10250 = frame (4k)
frame_vm_group_bin_10251 = frame (4k)
frame_vm_group_bin_10252 = frame (4k)
frame_vm_group_bin_10253 = frame (4k)
frame_vm_group_bin_10254 = frame (4k)
frame_vm_group_bin_10255 = frame (4k)
frame_vm_group_bin_10256 = frame (4k)
frame_vm_group_bin_10257 = frame (4k)
frame_vm_group_bin_10258 = frame (4k)
frame_vm_group_bin_10259 = frame (4k)
frame_vm_group_bin_1026 = frame (4k)
frame_vm_group_bin_10260 = frame (4k)
frame_vm_group_bin_10261 = frame (4k)
frame_vm_group_bin_10262 = frame (4k)
frame_vm_group_bin_10263 = frame (4k)
frame_vm_group_bin_10264 = frame (4k)
frame_vm_group_bin_10265 = frame (4k)
frame_vm_group_bin_10266 = frame (4k)
frame_vm_group_bin_10267 = frame (4k)
frame_vm_group_bin_10268 = frame (4k)
frame_vm_group_bin_10269 = frame (4k)
frame_vm_group_bin_1027 = frame (4k)
frame_vm_group_bin_10270 = frame (4k)
frame_vm_group_bin_10271 = frame (4k)
frame_vm_group_bin_10272 = frame (4k)
frame_vm_group_bin_10273 = frame (4k)
frame_vm_group_bin_10274 = frame (4k)
frame_vm_group_bin_10275 = frame (4k)
frame_vm_group_bin_10276 = frame (4k)
frame_vm_group_bin_10277 = frame (4k)
frame_vm_group_bin_10278 = frame (4k)
frame_vm_group_bin_10279 = frame (4k)
frame_vm_group_bin_1028 = frame (4k)
frame_vm_group_bin_10280 = frame (4k)
frame_vm_group_bin_10281 = frame (4k)
frame_vm_group_bin_10282 = frame (4k)
frame_vm_group_bin_10283 = frame (4k)
frame_vm_group_bin_10284 = frame (4k)
frame_vm_group_bin_10285 = frame (4k)
frame_vm_group_bin_10286 = frame (4k)
frame_vm_group_bin_10287 = frame (4k)
frame_vm_group_bin_10288 = frame (4k)
frame_vm_group_bin_10289 = frame (4k)
frame_vm_group_bin_1029 = frame (4k)
frame_vm_group_bin_10290 = frame (4k)
frame_vm_group_bin_10291 = frame (4k)
frame_vm_group_bin_10292 = frame (4k)
frame_vm_group_bin_10293 = frame (4k)
frame_vm_group_bin_10294 = frame (4k)
frame_vm_group_bin_10295 = frame (4k)
frame_vm_group_bin_10296 = frame (4k)
frame_vm_group_bin_10297 = frame (4k)
frame_vm_group_bin_10298 = frame (4k)
frame_vm_group_bin_10299 = frame (4k)
frame_vm_group_bin_1030 = frame (4k)
frame_vm_group_bin_10300 = frame (4k)
frame_vm_group_bin_10301 = frame (4k)
frame_vm_group_bin_10302 = frame (4k)
frame_vm_group_bin_10303 = frame (4k)
frame_vm_group_bin_10304 = frame (4k)
frame_vm_group_bin_10305 = frame (4k)
frame_vm_group_bin_10306 = frame (4k)
frame_vm_group_bin_10307 = frame (4k)
frame_vm_group_bin_10308 = frame (4k)
frame_vm_group_bin_10309 = frame (4k)
frame_vm_group_bin_1031 = frame (4k)
frame_vm_group_bin_10310 = frame (4k)
frame_vm_group_bin_10311 = frame (4k)
frame_vm_group_bin_10312 = frame (4k)
frame_vm_group_bin_10313 = frame (4k)
frame_vm_group_bin_10314 = frame (4k)
frame_vm_group_bin_10315 = frame (4k)
frame_vm_group_bin_10316 = frame (4k)
frame_vm_group_bin_10317 = frame (4k)
frame_vm_group_bin_10318 = frame (4k)
frame_vm_group_bin_10319 = frame (4k)
frame_vm_group_bin_1032 = frame (4k)
frame_vm_group_bin_10320 = frame (4k)
frame_vm_group_bin_10321 = frame (4k)
frame_vm_group_bin_10322 = frame (4k)
frame_vm_group_bin_10323 = frame (4k)
frame_vm_group_bin_10324 = frame (4k)
frame_vm_group_bin_10325 = frame (4k)
frame_vm_group_bin_10326 = frame (4k)
frame_vm_group_bin_10327 = frame (4k)
frame_vm_group_bin_10328 = frame (4k)
frame_vm_group_bin_10329 = frame (4k)
frame_vm_group_bin_1033 = frame (4k)
frame_vm_group_bin_10330 = frame (4k)
frame_vm_group_bin_10331 = frame (4k)
frame_vm_group_bin_10332 = frame (4k)
frame_vm_group_bin_10333 = frame (4k)
frame_vm_group_bin_10334 = frame (4k)
frame_vm_group_bin_10335 = frame (4k)
frame_vm_group_bin_10336 = frame (4k)
frame_vm_group_bin_10337 = frame (4k)
frame_vm_group_bin_10338 = frame (4k)
frame_vm_group_bin_10339 = frame (4k)
frame_vm_group_bin_1034 = frame (4k)
frame_vm_group_bin_10340 = frame (4k)
frame_vm_group_bin_10341 = frame (4k)
frame_vm_group_bin_10342 = frame (4k)
frame_vm_group_bin_10343 = frame (4k)
frame_vm_group_bin_10344 = frame (4k)
frame_vm_group_bin_10345 = frame (4k)
frame_vm_group_bin_10346 = frame (4k)
frame_vm_group_bin_10347 = frame (4k)
frame_vm_group_bin_10348 = frame (4k)
frame_vm_group_bin_10349 = frame (4k)
frame_vm_group_bin_1035 = frame (4k)
frame_vm_group_bin_10350 = frame (4k)
frame_vm_group_bin_10351 = frame (4k)
frame_vm_group_bin_10352 = frame (4k)
frame_vm_group_bin_10353 = frame (4k)
frame_vm_group_bin_10354 = frame (4k)
frame_vm_group_bin_10355 = frame (4k)
frame_vm_group_bin_10356 = frame (4k)
frame_vm_group_bin_10357 = frame (4k)
frame_vm_group_bin_10358 = frame (4k)
frame_vm_group_bin_10359 = frame (4k)
frame_vm_group_bin_1036 = frame (4k)
frame_vm_group_bin_10360 = frame (4k)
frame_vm_group_bin_10361 = frame (4k)
frame_vm_group_bin_10362 = frame (4k)
frame_vm_group_bin_10363 = frame (4k)
frame_vm_group_bin_10364 = frame (4k)
frame_vm_group_bin_10365 = frame (4k)
frame_vm_group_bin_10366 = frame (4k)
frame_vm_group_bin_10367 = frame (4k)
frame_vm_group_bin_10368 = frame (4k)
frame_vm_group_bin_10369 = frame (4k)
frame_vm_group_bin_1037 = frame (4k)
frame_vm_group_bin_10370 = frame (4k)
frame_vm_group_bin_10371 = frame (4k)
frame_vm_group_bin_10372 = frame (4k)
frame_vm_group_bin_10373 = frame (4k)
frame_vm_group_bin_10374 = frame (4k)
frame_vm_group_bin_10375 = frame (4k)
frame_vm_group_bin_10376 = frame (4k)
frame_vm_group_bin_10377 = frame (4k)
frame_vm_group_bin_10378 = frame (4k)
frame_vm_group_bin_10379 = frame (4k)
frame_vm_group_bin_1038 = frame (4k)
frame_vm_group_bin_10380 = frame (4k)
frame_vm_group_bin_10381 = frame (4k)
frame_vm_group_bin_10382 = frame (4k)
frame_vm_group_bin_10383 = frame (4k)
frame_vm_group_bin_10384 = frame (4k)
frame_vm_group_bin_10385 = frame (4k)
frame_vm_group_bin_10386 = frame (4k)
frame_vm_group_bin_10387 = frame (4k)
frame_vm_group_bin_10388 = frame (4k)
frame_vm_group_bin_10389 = frame (4k)
frame_vm_group_bin_1039 = frame (4k)
frame_vm_group_bin_10390 = frame (4k)
frame_vm_group_bin_10391 = frame (4k)
frame_vm_group_bin_10392 = frame (4k)
frame_vm_group_bin_10393 = frame (4k)
frame_vm_group_bin_10394 = frame (4k)
frame_vm_group_bin_10395 = frame (4k)
frame_vm_group_bin_10396 = frame (4k)
frame_vm_group_bin_10397 = frame (4k)
frame_vm_group_bin_10398 = frame (4k)
frame_vm_group_bin_10399 = frame (4k)
frame_vm_group_bin_1040 = frame (4k)
frame_vm_group_bin_10400 = frame (4k)
frame_vm_group_bin_10401 = frame (4k)
frame_vm_group_bin_10402 = frame (4k)
frame_vm_group_bin_10403 = frame (4k)
frame_vm_group_bin_10404 = frame (4k)
frame_vm_group_bin_10405 = frame (4k)
frame_vm_group_bin_10406 = frame (4k)
frame_vm_group_bin_10407 = frame (4k)
frame_vm_group_bin_10408 = frame (4k)
frame_vm_group_bin_10409 = frame (4k)
frame_vm_group_bin_1041 = frame (4k)
frame_vm_group_bin_10410 = frame (4k)
frame_vm_group_bin_10411 = frame (4k)
frame_vm_group_bin_10412 = frame (4k)
frame_vm_group_bin_10413 = frame (4k)
frame_vm_group_bin_10414 = frame (4k)
frame_vm_group_bin_10415 = frame (4k)
frame_vm_group_bin_10416 = frame (4k)
frame_vm_group_bin_10417 = frame (4k)
frame_vm_group_bin_10418 = frame (4k)
frame_vm_group_bin_10419 = frame (4k)
frame_vm_group_bin_1042 = frame (4k)
frame_vm_group_bin_10420 = frame (4k)
frame_vm_group_bin_10421 = frame (4k)
frame_vm_group_bin_10422 = frame (4k)
frame_vm_group_bin_10423 = frame (4k)
frame_vm_group_bin_10424 = frame (4k)
frame_vm_group_bin_10425 = frame (4k)
frame_vm_group_bin_10426 = frame (4k)
frame_vm_group_bin_10427 = frame (4k)
frame_vm_group_bin_10428 = frame (4k)
frame_vm_group_bin_10429 = frame (4k)
frame_vm_group_bin_1043 = frame (4k)
frame_vm_group_bin_10430 = frame (4k)
frame_vm_group_bin_10431 = frame (4k)
frame_vm_group_bin_10432 = frame (4k)
frame_vm_group_bin_10433 = frame (4k)
frame_vm_group_bin_10434 = frame (4k)
frame_vm_group_bin_10435 = frame (4k)
frame_vm_group_bin_10436 = frame (4k)
frame_vm_group_bin_10437 = frame (4k)
frame_vm_group_bin_10438 = frame (4k)
frame_vm_group_bin_10439 = frame (4k)
frame_vm_group_bin_1044 = frame (4k)
frame_vm_group_bin_10440 = frame (4k)
frame_vm_group_bin_10441 = frame (4k)
frame_vm_group_bin_10442 = frame (4k)
frame_vm_group_bin_10443 = frame (4k)
frame_vm_group_bin_10444 = frame (4k)
frame_vm_group_bin_10445 = frame (4k)
frame_vm_group_bin_10446 = frame (4k)
frame_vm_group_bin_10447 = frame (4k)
frame_vm_group_bin_10448 = frame (4k)
frame_vm_group_bin_10449 = frame (4k)
frame_vm_group_bin_1045 = frame (4k)
frame_vm_group_bin_10450 = frame (4k)
frame_vm_group_bin_10451 = frame (4k)
frame_vm_group_bin_10452 = frame (4k)
frame_vm_group_bin_10453 = frame (4k)
frame_vm_group_bin_10454 = frame (4k)
frame_vm_group_bin_10455 = frame (4k)
frame_vm_group_bin_10456 = frame (4k)
frame_vm_group_bin_10457 = frame (4k)
frame_vm_group_bin_10458 = frame (4k)
frame_vm_group_bin_10459 = frame (4k)
frame_vm_group_bin_1046 = frame (4k)
frame_vm_group_bin_10460 = frame (4k)
frame_vm_group_bin_10461 = frame (4k)
frame_vm_group_bin_10462 = frame (4k)
frame_vm_group_bin_10463 = frame (4k)
frame_vm_group_bin_10464 = frame (4k)
frame_vm_group_bin_10465 = frame (4k)
frame_vm_group_bin_10466 = frame (4k)
frame_vm_group_bin_10467 = frame (4k)
frame_vm_group_bin_10468 = frame (4k)
frame_vm_group_bin_10469 = frame (4k)
frame_vm_group_bin_1047 = frame (4k)
frame_vm_group_bin_10470 = frame (4k)
frame_vm_group_bin_10471 = frame (4k)
frame_vm_group_bin_10472 = frame (4k)
frame_vm_group_bin_10473 = frame (4k)
frame_vm_group_bin_10474 = frame (4k)
frame_vm_group_bin_10475 = frame (4k)
frame_vm_group_bin_10476 = frame (4k)
frame_vm_group_bin_10477 = frame (4k)
frame_vm_group_bin_10478 = frame (4k)
frame_vm_group_bin_10479 = frame (4k)
frame_vm_group_bin_1048 = frame (4k)
frame_vm_group_bin_10480 = frame (4k)
frame_vm_group_bin_10481 = frame (4k)
frame_vm_group_bin_10482 = frame (4k)
frame_vm_group_bin_10483 = frame (4k)
frame_vm_group_bin_10484 = frame (4k)
frame_vm_group_bin_10485 = frame (4k)
frame_vm_group_bin_10486 = frame (4k)
frame_vm_group_bin_10487 = frame (4k)
frame_vm_group_bin_10488 = frame (4k)
frame_vm_group_bin_10489 = frame (4k)
frame_vm_group_bin_1049 = frame (4k)
frame_vm_group_bin_10490 = frame (4k)
frame_vm_group_bin_10491 = frame (4k)
frame_vm_group_bin_10492 = frame (4k)
frame_vm_group_bin_10493 = frame (4k)
frame_vm_group_bin_10494 = frame (4k)
frame_vm_group_bin_10495 = frame (4k)
frame_vm_group_bin_10496 = frame (4k)
frame_vm_group_bin_10497 = frame (4k)
frame_vm_group_bin_10498 = frame (4k)
frame_vm_group_bin_10499 = frame (4k)
frame_vm_group_bin_1050 = frame (4k)
frame_vm_group_bin_10500 = frame (4k)
frame_vm_group_bin_10501 = frame (4k)
frame_vm_group_bin_10502 = frame (4k)
frame_vm_group_bin_10503 = frame (4k)
frame_vm_group_bin_10504 = frame (4k)
frame_vm_group_bin_10505 = frame (4k)
frame_vm_group_bin_10506 = frame (4k)
frame_vm_group_bin_10507 = frame (4k)
frame_vm_group_bin_10508 = frame (4k)
frame_vm_group_bin_10509 = frame (4k)
frame_vm_group_bin_1051 = frame (4k)
frame_vm_group_bin_10510 = frame (4k)
frame_vm_group_bin_10511 = frame (4k)
frame_vm_group_bin_10512 = frame (4k)
frame_vm_group_bin_10513 = frame (4k)
frame_vm_group_bin_10514 = frame (4k)
frame_vm_group_bin_10515 = frame (4k)
frame_vm_group_bin_10516 = frame (4k)
frame_vm_group_bin_10517 = frame (4k)
frame_vm_group_bin_10518 = frame (4k)
frame_vm_group_bin_10519 = frame (4k)
frame_vm_group_bin_1052 = frame (4k)
frame_vm_group_bin_10520 = frame (4k)
frame_vm_group_bin_10521 = frame (4k)
frame_vm_group_bin_10522 = frame (4k)
frame_vm_group_bin_10523 = frame (4k)
frame_vm_group_bin_10524 = frame (4k)
frame_vm_group_bin_10525 = frame (4k)
frame_vm_group_bin_10526 = frame (4k)
frame_vm_group_bin_10527 = frame (4k)
frame_vm_group_bin_10528 = frame (4k)
frame_vm_group_bin_10529 = frame (4k)
frame_vm_group_bin_1053 = frame (4k)
frame_vm_group_bin_10530 = frame (4k)
frame_vm_group_bin_10531 = frame (4k)
frame_vm_group_bin_10532 = frame (4k)
frame_vm_group_bin_10533 = frame (4k)
frame_vm_group_bin_10534 = frame (4k)
frame_vm_group_bin_10535 = frame (4k)
frame_vm_group_bin_10536 = frame (4k)
frame_vm_group_bin_10537 = frame (4k)
frame_vm_group_bin_10538 = frame (4k)
frame_vm_group_bin_10539 = frame (4k)
frame_vm_group_bin_1054 = frame (4k)
frame_vm_group_bin_10540 = frame (4k)
frame_vm_group_bin_10541 = frame (4k)
frame_vm_group_bin_10542 = frame (4k)
frame_vm_group_bin_10543 = frame (4k)
frame_vm_group_bin_10544 = frame (4k)
frame_vm_group_bin_10545 = frame (4k)
frame_vm_group_bin_10546 = frame (4k)
frame_vm_group_bin_10547 = frame (4k)
frame_vm_group_bin_10548 = frame (4k)
frame_vm_group_bin_10549 = frame (4k)
frame_vm_group_bin_1055 = frame (4k)
frame_vm_group_bin_10550 = frame (4k)
frame_vm_group_bin_10551 = frame (4k)
frame_vm_group_bin_10552 = frame (4k)
frame_vm_group_bin_10553 = frame (4k)
frame_vm_group_bin_10554 = frame (4k)
frame_vm_group_bin_10555 = frame (4k)
frame_vm_group_bin_10556 = frame (4k)
frame_vm_group_bin_10557 = frame (4k)
frame_vm_group_bin_10558 = frame (4k)
frame_vm_group_bin_10559 = frame (4k)
frame_vm_group_bin_1056 = frame (4k)
frame_vm_group_bin_10560 = frame (4k)
frame_vm_group_bin_10561 = frame (4k)
frame_vm_group_bin_10562 = frame (4k)
frame_vm_group_bin_10563 = frame (4k)
frame_vm_group_bin_10564 = frame (4k)
frame_vm_group_bin_10565 = frame (4k)
frame_vm_group_bin_10566 = frame (4k)
frame_vm_group_bin_10567 = frame (4k)
frame_vm_group_bin_10568 = frame (4k)
frame_vm_group_bin_10569 = frame (4k)
frame_vm_group_bin_1057 = frame (4k)
frame_vm_group_bin_10570 = frame (4k)
frame_vm_group_bin_10571 = frame (4k)
frame_vm_group_bin_10572 = frame (4k)
frame_vm_group_bin_10573 = frame (4k)
frame_vm_group_bin_10574 = frame (4k)
frame_vm_group_bin_10575 = frame (4k)
frame_vm_group_bin_10576 = frame (4k)
frame_vm_group_bin_10577 = frame (4k)
frame_vm_group_bin_10578 = frame (4k)
frame_vm_group_bin_10579 = frame (4k)
frame_vm_group_bin_1058 = frame (4k)
frame_vm_group_bin_10580 = frame (4k)
frame_vm_group_bin_10581 = frame (4k)
frame_vm_group_bin_10582 = frame (4k)
frame_vm_group_bin_10583 = frame (4k)
frame_vm_group_bin_10584 = frame (4k)
frame_vm_group_bin_10585 = frame (4k)
frame_vm_group_bin_10586 = frame (4k)
frame_vm_group_bin_10587 = frame (4k)
frame_vm_group_bin_10588 = frame (4k)
frame_vm_group_bin_10589 = frame (4k)
frame_vm_group_bin_1059 = frame (4k)
frame_vm_group_bin_10590 = frame (4k)
frame_vm_group_bin_10591 = frame (4k)
frame_vm_group_bin_10592 = frame (4k)
frame_vm_group_bin_10593 = frame (4k)
frame_vm_group_bin_10594 = frame (4k)
frame_vm_group_bin_10595 = frame (4k)
frame_vm_group_bin_10596 = frame (4k)
frame_vm_group_bin_10597 = frame (4k)
frame_vm_group_bin_10598 = frame (4k)
frame_vm_group_bin_10599 = frame (4k)
frame_vm_group_bin_1060 = frame (4k)
frame_vm_group_bin_10600 = frame (4k)
frame_vm_group_bin_10601 = frame (4k)
frame_vm_group_bin_10602 = frame (4k)
frame_vm_group_bin_10603 = frame (4k)
frame_vm_group_bin_10604 = frame (4k)
frame_vm_group_bin_10605 = frame (4k)
frame_vm_group_bin_10606 = frame (4k)
frame_vm_group_bin_10607 = frame (4k)
frame_vm_group_bin_10608 = frame (4k)
frame_vm_group_bin_10609 = frame (4k)
frame_vm_group_bin_1061 = frame (4k)
frame_vm_group_bin_10610 = frame (4k)
frame_vm_group_bin_10611 = frame (4k)
frame_vm_group_bin_10612 = frame (4k)
frame_vm_group_bin_10613 = frame (4k)
frame_vm_group_bin_10614 = frame (4k)
frame_vm_group_bin_10615 = frame (4k)
frame_vm_group_bin_10616 = frame (4k)
frame_vm_group_bin_10617 = frame (4k)
frame_vm_group_bin_10618 = frame (4k)
frame_vm_group_bin_10619 = frame (4k)
frame_vm_group_bin_1062 = frame (4k)
frame_vm_group_bin_10620 = frame (4k)
frame_vm_group_bin_10621 = frame (4k)
frame_vm_group_bin_10622 = frame (4k)
frame_vm_group_bin_10623 = frame (4k)
frame_vm_group_bin_10624 = frame (4k)
frame_vm_group_bin_10625 = frame (4k)
frame_vm_group_bin_10626 = frame (4k)
frame_vm_group_bin_10627 = frame (4k)
frame_vm_group_bin_10628 = frame (4k)
frame_vm_group_bin_10629 = frame (4k)
frame_vm_group_bin_1063 = frame (4k)
frame_vm_group_bin_10630 = frame (4k)
frame_vm_group_bin_10631 = frame (4k)
frame_vm_group_bin_10632 = frame (4k)
frame_vm_group_bin_10633 = frame (4k)
frame_vm_group_bin_10634 = frame (4k)
frame_vm_group_bin_10635 = frame (4k)
frame_vm_group_bin_10636 = frame (4k)
frame_vm_group_bin_10637 = frame (4k)
frame_vm_group_bin_10638 = frame (4k)
frame_vm_group_bin_10639 = frame (4k)
frame_vm_group_bin_1064 = frame (4k)
frame_vm_group_bin_10640 = frame (4k)
frame_vm_group_bin_10641 = frame (4k)
frame_vm_group_bin_10642 = frame (4k)
frame_vm_group_bin_10643 = frame (4k)
frame_vm_group_bin_10644 = frame (4k)
frame_vm_group_bin_10645 = frame (4k)
frame_vm_group_bin_10646 = frame (4k)
frame_vm_group_bin_10647 = frame (4k)
frame_vm_group_bin_10648 = frame (4k)
frame_vm_group_bin_10649 = frame (4k)
frame_vm_group_bin_1065 = frame (4k)
frame_vm_group_bin_10650 = frame (4k)
frame_vm_group_bin_10651 = frame (4k)
frame_vm_group_bin_10652 = frame (4k)
frame_vm_group_bin_10653 = frame (4k)
frame_vm_group_bin_10654 = frame (4k)
frame_vm_group_bin_10655 = frame (4k)
frame_vm_group_bin_10656 = frame (4k)
frame_vm_group_bin_10657 = frame (4k)
frame_vm_group_bin_10658 = frame (4k)
frame_vm_group_bin_10659 = frame (4k)
frame_vm_group_bin_1066 = frame (4k)
frame_vm_group_bin_10660 = frame (4k)
frame_vm_group_bin_10661 = frame (4k)
frame_vm_group_bin_10662 = frame (4k)
frame_vm_group_bin_10663 = frame (4k)
frame_vm_group_bin_10664 = frame (4k)
frame_vm_group_bin_10665 = frame (4k)
frame_vm_group_bin_10666 = frame (4k)
frame_vm_group_bin_10667 = frame (4k)
frame_vm_group_bin_10668 = frame (4k)
frame_vm_group_bin_10669 = frame (4k)
frame_vm_group_bin_1067 = frame (4k)
frame_vm_group_bin_10670 = frame (4k)
frame_vm_group_bin_10671 = frame (4k)
frame_vm_group_bin_10672 = frame (4k)
frame_vm_group_bin_10673 = frame (4k)
frame_vm_group_bin_10674 = frame (4k)
frame_vm_group_bin_10675 = frame (4k)
frame_vm_group_bin_10676 = frame (4k)
frame_vm_group_bin_10677 = frame (4k)
frame_vm_group_bin_10678 = frame (4k)
frame_vm_group_bin_10679 = frame (4k)
frame_vm_group_bin_1068 = frame (4k)
frame_vm_group_bin_10680 = frame (4k)
frame_vm_group_bin_10681 = frame (4k)
frame_vm_group_bin_10682 = frame (4k)
frame_vm_group_bin_10683 = frame (4k)
frame_vm_group_bin_10684 = frame (4k)
frame_vm_group_bin_10685 = frame (4k)
frame_vm_group_bin_10686 = frame (4k)
frame_vm_group_bin_10687 = frame (4k)
frame_vm_group_bin_10688 = frame (4k)
frame_vm_group_bin_10689 = frame (4k)
frame_vm_group_bin_1069 = frame (4k)
frame_vm_group_bin_10690 = frame (4k)
frame_vm_group_bin_10691 = frame (4k)
frame_vm_group_bin_10692 = frame (4k)
frame_vm_group_bin_10693 = frame (4k)
frame_vm_group_bin_10694 = frame (4k)
frame_vm_group_bin_10695 = frame (4k)
frame_vm_group_bin_10696 = frame (4k)
frame_vm_group_bin_10697 = frame (4k)
frame_vm_group_bin_10698 = frame (4k)
frame_vm_group_bin_10699 = frame (4k)
frame_vm_group_bin_1070 = frame (4k)
frame_vm_group_bin_10700 = frame (4k)
frame_vm_group_bin_10701 = frame (4k)
frame_vm_group_bin_10702 = frame (4k)
frame_vm_group_bin_10703 = frame (4k)
frame_vm_group_bin_10704 = frame (4k)
frame_vm_group_bin_10705 = frame (4k)
frame_vm_group_bin_10706 = frame (4k)
frame_vm_group_bin_10707 = frame (4k)
frame_vm_group_bin_10708 = frame (4k)
frame_vm_group_bin_10709 = frame (4k)
frame_vm_group_bin_1071 = frame (4k)
frame_vm_group_bin_10710 = frame (4k)
frame_vm_group_bin_10711 = frame (4k)
frame_vm_group_bin_10712 = frame (4k)
frame_vm_group_bin_10713 = frame (4k)
frame_vm_group_bin_10714 = frame (4k)
frame_vm_group_bin_10715 = frame (4k)
frame_vm_group_bin_10716 = frame (4k)
frame_vm_group_bin_10717 = frame (4k)
frame_vm_group_bin_10718 = frame (4k)
frame_vm_group_bin_10719 = frame (4k)
frame_vm_group_bin_1072 = frame (4k)
frame_vm_group_bin_10720 = frame (4k)
frame_vm_group_bin_10721 = frame (4k)
frame_vm_group_bin_10722 = frame (4k)
frame_vm_group_bin_10723 = frame (4k)
frame_vm_group_bin_10724 = frame (4k)
frame_vm_group_bin_10725 = frame (4k)
frame_vm_group_bin_10726 = frame (4k)
frame_vm_group_bin_10727 = frame (4k)
frame_vm_group_bin_10728 = frame (4k)
frame_vm_group_bin_10729 = frame (4k)
frame_vm_group_bin_1073 = frame (4k)
frame_vm_group_bin_10730 = frame (4k)
frame_vm_group_bin_10731 = frame (4k)
frame_vm_group_bin_10732 = frame (4k)
frame_vm_group_bin_10733 = frame (4k)
frame_vm_group_bin_10734 = frame (4k)
frame_vm_group_bin_10735 = frame (4k)
frame_vm_group_bin_10736 = frame (4k)
frame_vm_group_bin_10737 = frame (4k)
frame_vm_group_bin_10738 = frame (4k)
frame_vm_group_bin_10739 = frame (4k)
frame_vm_group_bin_1074 = frame (4k)
frame_vm_group_bin_10740 = frame (4k)
frame_vm_group_bin_10741 = frame (4k)
frame_vm_group_bin_10742 = frame (4k)
frame_vm_group_bin_10743 = frame (4k)
frame_vm_group_bin_10744 = frame (4k)
frame_vm_group_bin_10745 = frame (4k)
frame_vm_group_bin_10746 = frame (4k)
frame_vm_group_bin_10747 = frame (4k)
frame_vm_group_bin_10748 = frame (4k)
frame_vm_group_bin_10749 = frame (4k)
frame_vm_group_bin_1075 = frame (4k)
frame_vm_group_bin_10750 = frame (4k)
frame_vm_group_bin_10751 = frame (4k)
frame_vm_group_bin_10752 = frame (4k)
frame_vm_group_bin_10753 = frame (4k)
frame_vm_group_bin_10754 = frame (4k)
frame_vm_group_bin_10755 = frame (4k)
frame_vm_group_bin_10756 = frame (4k)
frame_vm_group_bin_10757 = frame (4k)
frame_vm_group_bin_10758 = frame (4k)
frame_vm_group_bin_10759 = frame (4k)
frame_vm_group_bin_1076 = frame (4k)
frame_vm_group_bin_10760 = frame (4k)
frame_vm_group_bin_10761 = frame (4k)
frame_vm_group_bin_10762 = frame (4k)
frame_vm_group_bin_10763 = frame (4k)
frame_vm_group_bin_10764 = frame (4k)
frame_vm_group_bin_10765 = frame (4k)
frame_vm_group_bin_10766 = frame (4k)
frame_vm_group_bin_10767 = frame (4k)
frame_vm_group_bin_10768 = frame (4k)
frame_vm_group_bin_10769 = frame (4k)
frame_vm_group_bin_1077 = frame (4k)
frame_vm_group_bin_10770 = frame (4k)
frame_vm_group_bin_10771 = frame (4k)
frame_vm_group_bin_10772 = frame (4k)
frame_vm_group_bin_10773 = frame (4k)
frame_vm_group_bin_10774 = frame (4k)
frame_vm_group_bin_10775 = frame (4k)
frame_vm_group_bin_10776 = frame (4k)
frame_vm_group_bin_10777 = frame (4k)
frame_vm_group_bin_10778 = frame (4k)
frame_vm_group_bin_10779 = frame (4k)
frame_vm_group_bin_1078 = frame (4k)
frame_vm_group_bin_10780 = frame (4k)
frame_vm_group_bin_10781 = frame (4k)
frame_vm_group_bin_10782 = frame (4k)
frame_vm_group_bin_10783 = frame (4k)
frame_vm_group_bin_10784 = frame (4k)
frame_vm_group_bin_10785 = frame (4k)
frame_vm_group_bin_10786 = frame (4k)
frame_vm_group_bin_10787 = frame (4k)
frame_vm_group_bin_10788 = frame (4k)
frame_vm_group_bin_10789 = frame (4k)
frame_vm_group_bin_1079 = frame (4k)
frame_vm_group_bin_10790 = frame (4k)
frame_vm_group_bin_10791 = frame (4k)
frame_vm_group_bin_10792 = frame (4k)
frame_vm_group_bin_10793 = frame (4k)
frame_vm_group_bin_10794 = frame (4k)
frame_vm_group_bin_10795 = frame (4k)
frame_vm_group_bin_10796 = frame (4k)
frame_vm_group_bin_10797 = frame (4k)
frame_vm_group_bin_10798 = frame (4k)
frame_vm_group_bin_10799 = frame (4k)
frame_vm_group_bin_1080 = frame (4k)
frame_vm_group_bin_10800 = frame (4k)
frame_vm_group_bin_10801 = frame (4k)
frame_vm_group_bin_10802 = frame (4k)
frame_vm_group_bin_10803 = frame (4k)
frame_vm_group_bin_10804 = frame (4k)
frame_vm_group_bin_10805 = frame (4k)
frame_vm_group_bin_10806 = frame (4k)
frame_vm_group_bin_10807 = frame (4k)
frame_vm_group_bin_10808 = frame (4k)
frame_vm_group_bin_10809 = frame (4k)
frame_vm_group_bin_1081 = frame (4k)
frame_vm_group_bin_10810 = frame (4k)
frame_vm_group_bin_10811 = frame (4k)
frame_vm_group_bin_10812 = frame (4k)
frame_vm_group_bin_10813 = frame (4k)
frame_vm_group_bin_10814 = frame (4k)
frame_vm_group_bin_10815 = frame (4k)
frame_vm_group_bin_10816 = frame (4k)
frame_vm_group_bin_10817 = frame (4k)
frame_vm_group_bin_10818 = frame (4k)
frame_vm_group_bin_10819 = frame (4k)
frame_vm_group_bin_1082 = frame (4k)
frame_vm_group_bin_10820 = frame (4k)
frame_vm_group_bin_10821 = frame (4k)
frame_vm_group_bin_10822 = frame (4k)
frame_vm_group_bin_10823 = frame (4k)
frame_vm_group_bin_10824 = frame (4k)
frame_vm_group_bin_10825 = frame (4k)
frame_vm_group_bin_10826 = frame (4k)
frame_vm_group_bin_10827 = frame (4k)
frame_vm_group_bin_10828 = frame (4k)
frame_vm_group_bin_10829 = frame (4k)
frame_vm_group_bin_1083 = frame (4k)
frame_vm_group_bin_10830 = frame (4k)
frame_vm_group_bin_10831 = frame (4k)
frame_vm_group_bin_10832 = frame (4k)
frame_vm_group_bin_10833 = frame (4k)
frame_vm_group_bin_10834 = frame (4k)
frame_vm_group_bin_10835 = frame (4k)
frame_vm_group_bin_10836 = frame (4k)
frame_vm_group_bin_10837 = frame (4k)
frame_vm_group_bin_10838 = frame (4k)
frame_vm_group_bin_10839 = frame (4k)
frame_vm_group_bin_1084 = frame (4k)
frame_vm_group_bin_10840 = frame (4k)
frame_vm_group_bin_10841 = frame (4k)
frame_vm_group_bin_10842 = frame (4k)
frame_vm_group_bin_10843 = frame (4k)
frame_vm_group_bin_10844 = frame (4k)
frame_vm_group_bin_10845 = frame (4k)
frame_vm_group_bin_10846 = frame (4k)
frame_vm_group_bin_10847 = frame (4k)
frame_vm_group_bin_10848 = frame (4k)
frame_vm_group_bin_10849 = frame (4k)
frame_vm_group_bin_1085 = frame (4k)
frame_vm_group_bin_10850 = frame (4k)
frame_vm_group_bin_10851 = frame (4k)
frame_vm_group_bin_10852 = frame (4k)
frame_vm_group_bin_10853 = frame (4k)
frame_vm_group_bin_10854 = frame (4k)
frame_vm_group_bin_10855 = frame (4k)
frame_vm_group_bin_10856 = frame (4k)
frame_vm_group_bin_10857 = frame (4k)
frame_vm_group_bin_10858 = frame (4k)
frame_vm_group_bin_10859 = frame (4k)
frame_vm_group_bin_1086 = frame (4k)
frame_vm_group_bin_10860 = frame (4k)
frame_vm_group_bin_10861 = frame (4k)
frame_vm_group_bin_10862 = frame (4k)
frame_vm_group_bin_10863 = frame (4k)
frame_vm_group_bin_10864 = frame (4k)
frame_vm_group_bin_10865 = frame (4k)
frame_vm_group_bin_10866 = frame (4k)
frame_vm_group_bin_10867 = frame (4k)
frame_vm_group_bin_10868 = frame (4k)
frame_vm_group_bin_10869 = frame (4k)
frame_vm_group_bin_1087 = frame (4k)
frame_vm_group_bin_10870 = frame (4k)
frame_vm_group_bin_10871 = frame (4k)
frame_vm_group_bin_10872 = frame (4k)
frame_vm_group_bin_10873 = frame (4k)
frame_vm_group_bin_10874 = frame (4k)
frame_vm_group_bin_10875 = frame (4k)
frame_vm_group_bin_10876 = frame (4k)
frame_vm_group_bin_10877 = frame (4k)
frame_vm_group_bin_10878 = frame (4k)
frame_vm_group_bin_10879 = frame (4k)
frame_vm_group_bin_1088 = frame (4k)
frame_vm_group_bin_10880 = frame (4k)
frame_vm_group_bin_10881 = frame (4k)
frame_vm_group_bin_10882 = frame (4k)
frame_vm_group_bin_10883 = frame (4k)
frame_vm_group_bin_10884 = frame (4k)
frame_vm_group_bin_10885 = frame (4k)
frame_vm_group_bin_10886 = frame (4k)
frame_vm_group_bin_10887 = frame (4k)
frame_vm_group_bin_10888 = frame (4k)
frame_vm_group_bin_10889 = frame (4k)
frame_vm_group_bin_1089 = frame (4k)
frame_vm_group_bin_10890 = frame (4k)
frame_vm_group_bin_10891 = frame (4k)
frame_vm_group_bin_10892 = frame (4k)
frame_vm_group_bin_10893 = frame (4k)
frame_vm_group_bin_10894 = frame (4k)
frame_vm_group_bin_10895 = frame (4k)
frame_vm_group_bin_10896 = frame (4k)
frame_vm_group_bin_10897 = frame (4k)
frame_vm_group_bin_10898 = frame (4k)
frame_vm_group_bin_10899 = frame (4k)
frame_vm_group_bin_1090 = frame (4k)
frame_vm_group_bin_10900 = frame (4k)
frame_vm_group_bin_10901 = frame (4k)
frame_vm_group_bin_10902 = frame (4k)
frame_vm_group_bin_10903 = frame (4k)
frame_vm_group_bin_10904 = frame (4k)
frame_vm_group_bin_10905 = frame (4k)
frame_vm_group_bin_10906 = frame (4k)
frame_vm_group_bin_10907 = frame (4k)
frame_vm_group_bin_10908 = frame (4k)
frame_vm_group_bin_10909 = frame (4k)
frame_vm_group_bin_1091 = frame (4k)
frame_vm_group_bin_10910 = frame (4k)
frame_vm_group_bin_10911 = frame (4k)
frame_vm_group_bin_10912 = frame (4k)
frame_vm_group_bin_10913 = frame (4k)
frame_vm_group_bin_10914 = frame (4k)
frame_vm_group_bin_10915 = frame (4k)
frame_vm_group_bin_10916 = frame (4k)
frame_vm_group_bin_10917 = frame (4k)
frame_vm_group_bin_10918 = frame (4k)
frame_vm_group_bin_10919 = frame (4k)
frame_vm_group_bin_1092 = frame (4k)
frame_vm_group_bin_10920 = frame (4k)
frame_vm_group_bin_10921 = frame (4k)
frame_vm_group_bin_10922 = frame (4k)
frame_vm_group_bin_10923 = frame (4k)
frame_vm_group_bin_10924 = frame (4k)
frame_vm_group_bin_10925 = frame (4k)
frame_vm_group_bin_10926 = frame (4k)
frame_vm_group_bin_10927 = frame (4k)
frame_vm_group_bin_10928 = frame (4k)
frame_vm_group_bin_10929 = frame (4k)
frame_vm_group_bin_1093 = frame (4k)
frame_vm_group_bin_10930 = frame (4k)
frame_vm_group_bin_10931 = frame (4k)
frame_vm_group_bin_10932 = frame (4k)
frame_vm_group_bin_10933 = frame (4k)
frame_vm_group_bin_10934 = frame (4k)
frame_vm_group_bin_10935 = frame (4k)
frame_vm_group_bin_10936 = frame (4k)
frame_vm_group_bin_10937 = frame (4k)
frame_vm_group_bin_10938 = frame (4k)
frame_vm_group_bin_10939 = frame (4k)
frame_vm_group_bin_1094 = frame (4k)
frame_vm_group_bin_10940 = frame (4k)
frame_vm_group_bin_10941 = frame (4k)
frame_vm_group_bin_10942 = frame (4k)
frame_vm_group_bin_10943 = frame (4k)
frame_vm_group_bin_10944 = frame (4k)
frame_vm_group_bin_10945 = frame (4k)
frame_vm_group_bin_10946 = frame (4k)
frame_vm_group_bin_10947 = frame (4k)
frame_vm_group_bin_10948 = frame (4k)
frame_vm_group_bin_10949 = frame (4k)
frame_vm_group_bin_1095 = frame (4k)
frame_vm_group_bin_10950 = frame (4k)
frame_vm_group_bin_10951 = frame (4k)
frame_vm_group_bin_10952 = frame (4k)
frame_vm_group_bin_10953 = frame (4k)
frame_vm_group_bin_10954 = frame (4k)
frame_vm_group_bin_10955 = frame (4k)
frame_vm_group_bin_10956 = frame (4k)
frame_vm_group_bin_10957 = frame (4k)
frame_vm_group_bin_10958 = frame (4k)
frame_vm_group_bin_10959 = frame (4k)
frame_vm_group_bin_1096 = frame (4k)
frame_vm_group_bin_10960 = frame (4k)
frame_vm_group_bin_10961 = frame (4k)
frame_vm_group_bin_10962 = frame (4k)
frame_vm_group_bin_10963 = frame (4k)
frame_vm_group_bin_10964 = frame (4k)
frame_vm_group_bin_10965 = frame (4k)
frame_vm_group_bin_10966 = frame (4k)
frame_vm_group_bin_10967 = frame (4k)
frame_vm_group_bin_10968 = frame (4k)
frame_vm_group_bin_10969 = frame (4k)
frame_vm_group_bin_1097 = frame (4k)
frame_vm_group_bin_10970 = frame (4k)
frame_vm_group_bin_10971 = frame (4k)
frame_vm_group_bin_10972 = frame (4k)
frame_vm_group_bin_10973 = frame (4k)
frame_vm_group_bin_10974 = frame (4k)
frame_vm_group_bin_10975 = frame (4k)
frame_vm_group_bin_10976 = frame (4k)
frame_vm_group_bin_10977 = frame (4k)
frame_vm_group_bin_10978 = frame (4k)
frame_vm_group_bin_10979 = frame (4k)
frame_vm_group_bin_1098 = frame (4k)
frame_vm_group_bin_10980 = frame (4k)
frame_vm_group_bin_10981 = frame (4k)
frame_vm_group_bin_10982 = frame (4k)
frame_vm_group_bin_10983 = frame (4k)
frame_vm_group_bin_10984 = frame (4k)
frame_vm_group_bin_10985 = frame (4k)
frame_vm_group_bin_10986 = frame (4k)
frame_vm_group_bin_10987 = frame (4k)
frame_vm_group_bin_10988 = frame (4k)
frame_vm_group_bin_10989 = frame (4k)
frame_vm_group_bin_1099 = frame (4k)
frame_vm_group_bin_10990 = frame (4k)
frame_vm_group_bin_10991 = frame (4k)
frame_vm_group_bin_10992 = frame (4k)
frame_vm_group_bin_10993 = frame (4k)
frame_vm_group_bin_10994 = frame (4k)
frame_vm_group_bin_10995 = frame (4k)
frame_vm_group_bin_10996 = frame (4k)
frame_vm_group_bin_10997 = frame (4k)
frame_vm_group_bin_10998 = frame (4k)
frame_vm_group_bin_10999 = frame (4k)
frame_vm_group_bin_1100 = frame (4k)
frame_vm_group_bin_11000 = frame (4k)
frame_vm_group_bin_11001 = frame (4k)
frame_vm_group_bin_11002 = frame (4k)
frame_vm_group_bin_11003 = frame (4k)
frame_vm_group_bin_11004 = frame (4k)
frame_vm_group_bin_11005 = frame (4k)
frame_vm_group_bin_11006 = frame (4k)
frame_vm_group_bin_11007 = frame (4k)
frame_vm_group_bin_11008 = frame (4k)
frame_vm_group_bin_11009 = frame (4k)
frame_vm_group_bin_1101 = frame (4k)
frame_vm_group_bin_11010 = frame (4k)
frame_vm_group_bin_11011 = frame (4k)
frame_vm_group_bin_11012 = frame (4k)
frame_vm_group_bin_11013 = frame (4k)
frame_vm_group_bin_11014 = frame (4k)
frame_vm_group_bin_11015 = frame (4k)
frame_vm_group_bin_11016 = frame (4k)
frame_vm_group_bin_11017 = frame (4k)
frame_vm_group_bin_11018 = frame (4k)
frame_vm_group_bin_11019 = frame (4k)
frame_vm_group_bin_1102 = frame (4k)
frame_vm_group_bin_11020 = frame (4k)
frame_vm_group_bin_11021 = frame (4k)
frame_vm_group_bin_11022 = frame (4k)
frame_vm_group_bin_11023 = frame (4k)
frame_vm_group_bin_11024 = frame (4k)
frame_vm_group_bin_11025 = frame (4k)
frame_vm_group_bin_11026 = frame (4k)
frame_vm_group_bin_11027 = frame (4k)
frame_vm_group_bin_11028 = frame (4k)
frame_vm_group_bin_11029 = frame (4k)
frame_vm_group_bin_1103 = frame (4k)
frame_vm_group_bin_11030 = frame (4k)
frame_vm_group_bin_11031 = frame (4k)
frame_vm_group_bin_11032 = frame (4k)
frame_vm_group_bin_11033 = frame (4k)
frame_vm_group_bin_11034 = frame (4k)
frame_vm_group_bin_11035 = frame (4k)
frame_vm_group_bin_11036 = frame (4k)
frame_vm_group_bin_11037 = frame (4k)
frame_vm_group_bin_11038 = frame (4k)
frame_vm_group_bin_11039 = frame (4k)
frame_vm_group_bin_1104 = frame (4k)
frame_vm_group_bin_11040 = frame (4k)
frame_vm_group_bin_11041 = frame (4k)
frame_vm_group_bin_11042 = frame (4k)
frame_vm_group_bin_11043 = frame (4k)
frame_vm_group_bin_11044 = frame (4k)
frame_vm_group_bin_11045 = frame (4k)
frame_vm_group_bin_11046 = frame (4k)
frame_vm_group_bin_11047 = frame (4k)
frame_vm_group_bin_11048 = frame (4k)
frame_vm_group_bin_11049 = frame (4k)
frame_vm_group_bin_1105 = frame (4k)
frame_vm_group_bin_11050 = frame (4k)
frame_vm_group_bin_11051 = frame (4k)
frame_vm_group_bin_11052 = frame (4k)
frame_vm_group_bin_11053 = frame (4k)
frame_vm_group_bin_11054 = frame (4k)
frame_vm_group_bin_11055 = frame (4k)
frame_vm_group_bin_11056 = frame (4k)
frame_vm_group_bin_11057 = frame (4k)
frame_vm_group_bin_11058 = frame (4k)
frame_vm_group_bin_11059 = frame (4k)
frame_vm_group_bin_1106 = frame (4k)
frame_vm_group_bin_11060 = frame (4k)
frame_vm_group_bin_11061 = frame (4k)
frame_vm_group_bin_11062 = frame (4k)
frame_vm_group_bin_11063 = frame (4k)
frame_vm_group_bin_11064 = frame (4k)
frame_vm_group_bin_11065 = frame (4k)
frame_vm_group_bin_11066 = frame (4k)
frame_vm_group_bin_11067 = frame (4k)
frame_vm_group_bin_11068 = frame (4k)
frame_vm_group_bin_11069 = frame (4k)
frame_vm_group_bin_1107 = frame (4k)
frame_vm_group_bin_11070 = frame (4k)
frame_vm_group_bin_11071 = frame (4k)
frame_vm_group_bin_11072 = frame (4k)
frame_vm_group_bin_11073 = frame (4k)
frame_vm_group_bin_11074 = frame (4k)
frame_vm_group_bin_11075 = frame (4k)
frame_vm_group_bin_11076 = frame (4k)
frame_vm_group_bin_11077 = frame (4k)
frame_vm_group_bin_11078 = frame (4k)
frame_vm_group_bin_11079 = frame (4k)
frame_vm_group_bin_1108 = frame (4k)
frame_vm_group_bin_11080 = frame (4k)
frame_vm_group_bin_11081 = frame (4k)
frame_vm_group_bin_11082 = frame (4k)
frame_vm_group_bin_11083 = frame (4k)
frame_vm_group_bin_11084 = frame (4k)
frame_vm_group_bin_11085 = frame (4k)
frame_vm_group_bin_11086 = frame (4k)
frame_vm_group_bin_11087 = frame (4k)
frame_vm_group_bin_11088 = frame (4k)
frame_vm_group_bin_11089 = frame (4k)
frame_vm_group_bin_1109 = frame (4k)
frame_vm_group_bin_11090 = frame (4k)
frame_vm_group_bin_11091 = frame (4k)
frame_vm_group_bin_11092 = frame (4k)
frame_vm_group_bin_11093 = frame (4k)
frame_vm_group_bin_11094 = frame (4k)
frame_vm_group_bin_11095 = frame (4k)
frame_vm_group_bin_11096 = frame (4k)
frame_vm_group_bin_11097 = frame (4k)
frame_vm_group_bin_11098 = frame (4k)
frame_vm_group_bin_11099 = frame (4k)
frame_vm_group_bin_1110 = frame (4k)
frame_vm_group_bin_11100 = frame (4k)
frame_vm_group_bin_11101 = frame (4k)
frame_vm_group_bin_11102 = frame (4k)
frame_vm_group_bin_11103 = frame (4k)
frame_vm_group_bin_11104 = frame (4k)
frame_vm_group_bin_11105 = frame (4k)
frame_vm_group_bin_11106 = frame (4k)
frame_vm_group_bin_11107 = frame (4k)
frame_vm_group_bin_11108 = frame (4k)
frame_vm_group_bin_11109 = frame (4k)
frame_vm_group_bin_1111 = frame (4k)
frame_vm_group_bin_11110 = frame (4k)
frame_vm_group_bin_11111 = frame (4k)
frame_vm_group_bin_11112 = frame (4k)
frame_vm_group_bin_11113 = frame (4k)
frame_vm_group_bin_11114 = frame (4k)
frame_vm_group_bin_11115 = frame (4k)
frame_vm_group_bin_11116 = frame (4k)
frame_vm_group_bin_11117 = frame (4k)
frame_vm_group_bin_11118 = frame (4k)
frame_vm_group_bin_11119 = frame (4k)
frame_vm_group_bin_1112 = frame (4k)
frame_vm_group_bin_11120 = frame (4k)
frame_vm_group_bin_11121 = frame (4k)
frame_vm_group_bin_11122 = frame (4k)
frame_vm_group_bin_11123 = frame (4k)
frame_vm_group_bin_11124 = frame (4k)
frame_vm_group_bin_11125 = frame (4k)
frame_vm_group_bin_11126 = frame (4k)
frame_vm_group_bin_11127 = frame (4k)
frame_vm_group_bin_11128 = frame (4k)
frame_vm_group_bin_11129 = frame (4k)
frame_vm_group_bin_1113 = frame (4k)
frame_vm_group_bin_11130 = frame (4k)
frame_vm_group_bin_11131 = frame (4k)
frame_vm_group_bin_11132 = frame (4k)
frame_vm_group_bin_11133 = frame (4k)
frame_vm_group_bin_11134 = frame (4k)
frame_vm_group_bin_11135 = frame (4k)
frame_vm_group_bin_11136 = frame (4k)
frame_vm_group_bin_11137 = frame (4k)
frame_vm_group_bin_11138 = frame (4k)
frame_vm_group_bin_11139 = frame (4k)
frame_vm_group_bin_1114 = frame (4k)
frame_vm_group_bin_11140 = frame (4k)
frame_vm_group_bin_11141 = frame (4k)
frame_vm_group_bin_11142 = frame (4k)
frame_vm_group_bin_11143 = frame (4k)
frame_vm_group_bin_11144 = frame (4k)
frame_vm_group_bin_11145 = frame (4k)
frame_vm_group_bin_11146 = frame (4k)
frame_vm_group_bin_11147 = frame (4k)
frame_vm_group_bin_11148 = frame (4k)
frame_vm_group_bin_11149 = frame (4k)
frame_vm_group_bin_1115 = frame (4k)
frame_vm_group_bin_11150 = frame (4k)
frame_vm_group_bin_11151 = frame (4k)
frame_vm_group_bin_11152 = frame (4k)
frame_vm_group_bin_11153 = frame (4k)
frame_vm_group_bin_11154 = frame (4k)
frame_vm_group_bin_11155 = frame (4k)
frame_vm_group_bin_11156 = frame (4k)
frame_vm_group_bin_11157 = frame (4k)
frame_vm_group_bin_11158 = frame (4k)
frame_vm_group_bin_11159 = frame (4k)
frame_vm_group_bin_1116 = frame (4k)
frame_vm_group_bin_11160 = frame (4k)
frame_vm_group_bin_11161 = frame (4k)
frame_vm_group_bin_11162 = frame (4k)
frame_vm_group_bin_11163 = frame (4k)
frame_vm_group_bin_11164 = frame (4k)
frame_vm_group_bin_11165 = frame (4k)
frame_vm_group_bin_11166 = frame (4k)
frame_vm_group_bin_11167 = frame (4k)
frame_vm_group_bin_11168 = frame (4k)
frame_vm_group_bin_11169 = frame (4k)
frame_vm_group_bin_1117 = frame (4k)
frame_vm_group_bin_11170 = frame (4k)
frame_vm_group_bin_11171 = frame (4k)
frame_vm_group_bin_11172 = frame (4k)
frame_vm_group_bin_11173 = frame (4k)
frame_vm_group_bin_11174 = frame (4k)
frame_vm_group_bin_11175 = frame (4k)
frame_vm_group_bin_11176 = frame (4k)
frame_vm_group_bin_11177 = frame (4k)
frame_vm_group_bin_11178 = frame (4k)
frame_vm_group_bin_11179 = frame (4k)
frame_vm_group_bin_1118 = frame (4k)
frame_vm_group_bin_11180 = frame (4k)
frame_vm_group_bin_11181 = frame (4k)
frame_vm_group_bin_11182 = frame (4k)
frame_vm_group_bin_11183 = frame (4k)
frame_vm_group_bin_11184 = frame (4k)
frame_vm_group_bin_11185 = frame (4k)
frame_vm_group_bin_11186 = frame (4k)
frame_vm_group_bin_11187 = frame (4k)
frame_vm_group_bin_11188 = frame (4k)
frame_vm_group_bin_11189 = frame (4k)
frame_vm_group_bin_1119 = frame (4k)
frame_vm_group_bin_11190 = frame (4k)
frame_vm_group_bin_11191 = frame (4k)
frame_vm_group_bin_11192 = frame (4k)
frame_vm_group_bin_11193 = frame (4k)
frame_vm_group_bin_11194 = frame (4k)
frame_vm_group_bin_11195 = frame (4k)
frame_vm_group_bin_11196 = frame (4k)
frame_vm_group_bin_11197 = frame (4k)
frame_vm_group_bin_11198 = frame (4k)
frame_vm_group_bin_11199 = frame (4k)
frame_vm_group_bin_1120 = frame (4k)
frame_vm_group_bin_11200 = frame (4k)
frame_vm_group_bin_11201 = frame (4k)
frame_vm_group_bin_11202 = frame (4k)
frame_vm_group_bin_11203 = frame (4k)
frame_vm_group_bin_11204 = frame (4k)
frame_vm_group_bin_11205 = frame (4k)
frame_vm_group_bin_11206 = frame (4k)
frame_vm_group_bin_11207 = frame (4k)
frame_vm_group_bin_11208 = frame (4k)
frame_vm_group_bin_11209 = frame (4k)
frame_vm_group_bin_1121 = frame (4k)
frame_vm_group_bin_11210 = frame (4k)
frame_vm_group_bin_11211 = frame (4k)
frame_vm_group_bin_11212 = frame (4k)
frame_vm_group_bin_11213 = frame (4k)
frame_vm_group_bin_11214 = frame (4k)
frame_vm_group_bin_11215 = frame (4k)
frame_vm_group_bin_11216 = frame (4k)
frame_vm_group_bin_11217 = frame (4k)
frame_vm_group_bin_11218 = frame (4k)
frame_vm_group_bin_11219 = frame (4k)
frame_vm_group_bin_1122 = frame (4k)
frame_vm_group_bin_11220 = frame (4k)
frame_vm_group_bin_11221 = frame (4k)
frame_vm_group_bin_11222 = frame (4k)
frame_vm_group_bin_11223 = frame (4k)
frame_vm_group_bin_11224 = frame (4k)
frame_vm_group_bin_11225 = frame (4k)
frame_vm_group_bin_11226 = frame (4k)
frame_vm_group_bin_11227 = frame (4k)
frame_vm_group_bin_11228 = frame (4k)
frame_vm_group_bin_11229 = frame (4k)
frame_vm_group_bin_1123 = frame (4k)
frame_vm_group_bin_11230 = frame (4k)
frame_vm_group_bin_11231 = frame (4k)
frame_vm_group_bin_11232 = frame (4k)
frame_vm_group_bin_11233 = frame (4k)
frame_vm_group_bin_11234 = frame (4k)
frame_vm_group_bin_11235 = frame (4k)
frame_vm_group_bin_11236 = frame (4k)
frame_vm_group_bin_11237 = frame (4k)
frame_vm_group_bin_11238 = frame (4k)
frame_vm_group_bin_11239 = frame (4k)
frame_vm_group_bin_1124 = frame (4k)
frame_vm_group_bin_11240 = frame (4k)
frame_vm_group_bin_11241 = frame (4k)
frame_vm_group_bin_11242 = frame (4k)
frame_vm_group_bin_11243 = frame (4k)
frame_vm_group_bin_11244 = frame (4k)
frame_vm_group_bin_11245 = frame (4k)
frame_vm_group_bin_11246 = frame (4k)
frame_vm_group_bin_11247 = frame (4k)
frame_vm_group_bin_11248 = frame (4k)
frame_vm_group_bin_11249 = frame (4k)
frame_vm_group_bin_1125 = frame (4k)
frame_vm_group_bin_11250 = frame (4k)
frame_vm_group_bin_11251 = frame (4k)
frame_vm_group_bin_11252 = frame (4k)
frame_vm_group_bin_11253 = frame (4k)
frame_vm_group_bin_11254 = frame (4k)
frame_vm_group_bin_11255 = frame (4k)
frame_vm_group_bin_11256 = frame (4k)
frame_vm_group_bin_11257 = frame (4k)
frame_vm_group_bin_11258 = frame (4k)
frame_vm_group_bin_11259 = frame (4k)
frame_vm_group_bin_1126 = frame (4k)
frame_vm_group_bin_11260 = frame (4k)
frame_vm_group_bin_11261 = frame (4k)
frame_vm_group_bin_11262 = frame (4k)
frame_vm_group_bin_11263 = frame (4k)
frame_vm_group_bin_11264 = frame (4k)
frame_vm_group_bin_11265 = frame (4k)
frame_vm_group_bin_11266 = frame (4k)
frame_vm_group_bin_11267 = frame (4k)
frame_vm_group_bin_11268 = frame (4k)
frame_vm_group_bin_11269 = frame (4k)
frame_vm_group_bin_1127 = frame (4k)
frame_vm_group_bin_11270 = frame (4k)
frame_vm_group_bin_11271 = frame (4k)
frame_vm_group_bin_11272 = frame (4k)
frame_vm_group_bin_11273 = frame (4k)
frame_vm_group_bin_11274 = frame (4k)
frame_vm_group_bin_11275 = frame (4k)
frame_vm_group_bin_11276 = frame (4k)
frame_vm_group_bin_11277 = frame (4k)
frame_vm_group_bin_11278 = frame (4k)
frame_vm_group_bin_11279 = frame (4k)
frame_vm_group_bin_1128 = frame (4k)
frame_vm_group_bin_11280 = frame (4k)
frame_vm_group_bin_11281 = frame (4k)
frame_vm_group_bin_11282 = frame (4k)
frame_vm_group_bin_11283 = frame (4k)
frame_vm_group_bin_11284 = frame (4k)
frame_vm_group_bin_11285 = frame (4k)
frame_vm_group_bin_11286 = frame (4k)
frame_vm_group_bin_11287 = frame (4k)
frame_vm_group_bin_11288 = frame (4k)
frame_vm_group_bin_11289 = frame (4k)
frame_vm_group_bin_1129 = frame (4k)
frame_vm_group_bin_11290 = frame (4k)
frame_vm_group_bin_11291 = frame (4k)
frame_vm_group_bin_11292 = frame (4k)
frame_vm_group_bin_11293 = frame (4k)
frame_vm_group_bin_11294 = frame (4k)
frame_vm_group_bin_11295 = frame (4k)
frame_vm_group_bin_11296 = frame (4k)
frame_vm_group_bin_11297 = frame (4k)
frame_vm_group_bin_11298 = frame (4k)
frame_vm_group_bin_11299 = frame (4k)
frame_vm_group_bin_1130 = frame (4k)
frame_vm_group_bin_11300 = frame (4k)
frame_vm_group_bin_11301 = frame (4k)
frame_vm_group_bin_11302 = frame (4k)
frame_vm_group_bin_11303 = frame (4k)
frame_vm_group_bin_11304 = frame (4k)
frame_vm_group_bin_11305 = frame (4k)
frame_vm_group_bin_11306 = frame (4k)
frame_vm_group_bin_11307 = frame (4k)
frame_vm_group_bin_11308 = frame (4k)
frame_vm_group_bin_11309 = frame (4k)
frame_vm_group_bin_1131 = frame (4k)
frame_vm_group_bin_11310 = frame (4k)
frame_vm_group_bin_11311 = frame (4k)
frame_vm_group_bin_11312 = frame (4k)
frame_vm_group_bin_11313 = frame (4k)
frame_vm_group_bin_11314 = frame (4k)
frame_vm_group_bin_11315 = frame (4k)
frame_vm_group_bin_11316 = frame (4k)
frame_vm_group_bin_11317 = frame (4k)
frame_vm_group_bin_11318 = frame (4k)
frame_vm_group_bin_11319 = frame (4k)
frame_vm_group_bin_1132 = frame (4k)
frame_vm_group_bin_11320 = frame (4k)
frame_vm_group_bin_11321 = frame (4k)
frame_vm_group_bin_11322 = frame (4k)
frame_vm_group_bin_11323 = frame (4k)
frame_vm_group_bin_11324 = frame (4k)
frame_vm_group_bin_11325 = frame (4k)
frame_vm_group_bin_11326 = frame (4k)
frame_vm_group_bin_11327 = frame (4k)
frame_vm_group_bin_11328 = frame (4k)
frame_vm_group_bin_11329 = frame (4k)
frame_vm_group_bin_1133 = frame (4k)
frame_vm_group_bin_11330 = frame (4k)
frame_vm_group_bin_11331 = frame (4k)
frame_vm_group_bin_11332 = frame (4k)
frame_vm_group_bin_11333 = frame (4k)
frame_vm_group_bin_11334 = frame (4k)
frame_vm_group_bin_11335 = frame (4k)
frame_vm_group_bin_11336 = frame (4k)
frame_vm_group_bin_11337 = frame (4k)
frame_vm_group_bin_11338 = frame (4k)
frame_vm_group_bin_11339 = frame (4k)
frame_vm_group_bin_1134 = frame (4k)
frame_vm_group_bin_11340 = frame (4k)
frame_vm_group_bin_11341 = frame (4k)
frame_vm_group_bin_11342 = frame (4k)
frame_vm_group_bin_11343 = frame (4k)
frame_vm_group_bin_11344 = frame (4k)
frame_vm_group_bin_11345 = frame (4k)
frame_vm_group_bin_11346 = frame (4k)
frame_vm_group_bin_11347 = frame (4k)
frame_vm_group_bin_11348 = frame (4k)
frame_vm_group_bin_11349 = frame (4k)
frame_vm_group_bin_1135 = frame (4k)
frame_vm_group_bin_11350 = frame (4k)
frame_vm_group_bin_11351 = frame (4k)
frame_vm_group_bin_11352 = frame (4k)
frame_vm_group_bin_11353 = frame (4k)
frame_vm_group_bin_11354 = frame (4k)
frame_vm_group_bin_11355 = frame (4k)
frame_vm_group_bin_11356 = frame (4k)
frame_vm_group_bin_11357 = frame (4k)
frame_vm_group_bin_11358 = frame (4k)
frame_vm_group_bin_11359 = frame (4k)
frame_vm_group_bin_1136 = frame (4k)
frame_vm_group_bin_11360 = frame (4k)
frame_vm_group_bin_11361 = frame (4k)
frame_vm_group_bin_11362 = frame (4k)
frame_vm_group_bin_11363 = frame (4k)
frame_vm_group_bin_11364 = frame (4k)
frame_vm_group_bin_11365 = frame (4k)
frame_vm_group_bin_11366 = frame (4k)
frame_vm_group_bin_11367 = frame (4k)
frame_vm_group_bin_11368 = frame (4k)
frame_vm_group_bin_11369 = frame (4k)
frame_vm_group_bin_1137 = frame (4k)
frame_vm_group_bin_11370 = frame (4k)
frame_vm_group_bin_11371 = frame (4k)
frame_vm_group_bin_11372 = frame (4k)
frame_vm_group_bin_11373 = frame (4k)
frame_vm_group_bin_11374 = frame (4k)
frame_vm_group_bin_11375 = frame (4k)
frame_vm_group_bin_11376 = frame (4k)
frame_vm_group_bin_11377 = frame (4k)
frame_vm_group_bin_11378 = frame (4k)
frame_vm_group_bin_11379 = frame (4k)
frame_vm_group_bin_1138 = frame (4k)
frame_vm_group_bin_11380 = frame (4k)
frame_vm_group_bin_11381 = frame (4k)
frame_vm_group_bin_11382 = frame (4k)
frame_vm_group_bin_11383 = frame (4k)
frame_vm_group_bin_11384 = frame (4k)
frame_vm_group_bin_11385 = frame (4k)
frame_vm_group_bin_11386 = frame (4k)
frame_vm_group_bin_11387 = frame (4k)
frame_vm_group_bin_11388 = frame (4k)
frame_vm_group_bin_11389 = frame (4k)
frame_vm_group_bin_1139 = frame (4k)
frame_vm_group_bin_11390 = frame (4k)
frame_vm_group_bin_11391 = frame (4k)
frame_vm_group_bin_11392 = frame (4k)
frame_vm_group_bin_11393 = frame (4k)
frame_vm_group_bin_11394 = frame (4k)
frame_vm_group_bin_11395 = frame (4k)
frame_vm_group_bin_11396 = frame (4k)
frame_vm_group_bin_11397 = frame (4k)
frame_vm_group_bin_11398 = frame (4k)
frame_vm_group_bin_11399 = frame (4k)
frame_vm_group_bin_1140 = frame (4k)
frame_vm_group_bin_11400 = frame (4k)
frame_vm_group_bin_11401 = frame (4k)
frame_vm_group_bin_11402 = frame (4k)
frame_vm_group_bin_11403 = frame (4k)
frame_vm_group_bin_11404 = frame (4k)
frame_vm_group_bin_11405 = frame (4k)
frame_vm_group_bin_11406 = frame (4k)
frame_vm_group_bin_11407 = frame (4k)
frame_vm_group_bin_11408 = frame (4k)
frame_vm_group_bin_11409 = frame (4k)
frame_vm_group_bin_1141 = frame (4k)
frame_vm_group_bin_11410 = frame (4k)
frame_vm_group_bin_11411 = frame (4k)
frame_vm_group_bin_11412 = frame (4k)
frame_vm_group_bin_11413 = frame (4k)
frame_vm_group_bin_11414 = frame (4k)
frame_vm_group_bin_11415 = frame (4k)
frame_vm_group_bin_11416 = frame (4k)
frame_vm_group_bin_11417 = frame (4k)
frame_vm_group_bin_11418 = frame (4k)
frame_vm_group_bin_11419 = frame (4k)
frame_vm_group_bin_1142 = frame (4k)
frame_vm_group_bin_11420 = frame (4k)
frame_vm_group_bin_11421 = frame (4k)
frame_vm_group_bin_11422 = frame (4k)
frame_vm_group_bin_11423 = frame (4k)
frame_vm_group_bin_11424 = frame (4k)
frame_vm_group_bin_11425 = frame (4k)
frame_vm_group_bin_11426 = frame (4k)
frame_vm_group_bin_11427 = frame (4k)
frame_vm_group_bin_11428 = frame (4k)
frame_vm_group_bin_11429 = frame (4k)
frame_vm_group_bin_1143 = frame (4k)
frame_vm_group_bin_11430 = frame (4k)
frame_vm_group_bin_11431 = frame (4k)
frame_vm_group_bin_11432 = frame (4k)
frame_vm_group_bin_11433 = frame (4k)
frame_vm_group_bin_11434 = frame (4k)
frame_vm_group_bin_11435 = frame (4k)
frame_vm_group_bin_11436 = frame (4k)
frame_vm_group_bin_11437 = frame (4k)
frame_vm_group_bin_11438 = frame (4k)
frame_vm_group_bin_11439 = frame (4k)
frame_vm_group_bin_1144 = frame (4k)
frame_vm_group_bin_11440 = frame (4k)
frame_vm_group_bin_11441 = frame (4k)
frame_vm_group_bin_11442 = frame (4k)
frame_vm_group_bin_11443 = frame (4k)
frame_vm_group_bin_11444 = frame (4k)
frame_vm_group_bin_11445 = frame (4k)
frame_vm_group_bin_11446 = frame (4k)
frame_vm_group_bin_11447 = frame (4k)
frame_vm_group_bin_11448 = frame (4k)
frame_vm_group_bin_11449 = frame (4k)
frame_vm_group_bin_1145 = frame (4k)
frame_vm_group_bin_11450 = frame (4k)
frame_vm_group_bin_11451 = frame (4k)
frame_vm_group_bin_11452 = frame (4k)
frame_vm_group_bin_11453 = frame (4k)
frame_vm_group_bin_11454 = frame (4k)
frame_vm_group_bin_11455 = frame (4k)
frame_vm_group_bin_11456 = frame (4k)
frame_vm_group_bin_11457 = frame (4k)
frame_vm_group_bin_11458 = frame (4k)
frame_vm_group_bin_11459 = frame (4k)
frame_vm_group_bin_1146 = frame (4k)
frame_vm_group_bin_11460 = frame (4k)
frame_vm_group_bin_11461 = frame (4k)
frame_vm_group_bin_11462 = frame (4k)
frame_vm_group_bin_11463 = frame (4k)
frame_vm_group_bin_11464 = frame (4k)
frame_vm_group_bin_11465 = frame (4k)
frame_vm_group_bin_11466 = frame (4k)
frame_vm_group_bin_11467 = frame (4k)
frame_vm_group_bin_11468 = frame (4k)
frame_vm_group_bin_11469 = frame (4k)
frame_vm_group_bin_1147 = frame (4k)
frame_vm_group_bin_11470 = frame (4k)
frame_vm_group_bin_11471 = frame (4k)
frame_vm_group_bin_11472 = frame (4k)
frame_vm_group_bin_11473 = frame (4k)
frame_vm_group_bin_11474 = frame (4k)
frame_vm_group_bin_11475 = frame (4k)
frame_vm_group_bin_11476 = frame (4k)
frame_vm_group_bin_11477 = frame (4k)
frame_vm_group_bin_11478 = frame (4k)
frame_vm_group_bin_11479 = frame (4k)
frame_vm_group_bin_1148 = frame (4k)
frame_vm_group_bin_11480 = frame (4k)
frame_vm_group_bin_11481 = frame (4k)
frame_vm_group_bin_11482 = frame (4k)
frame_vm_group_bin_11483 = frame (4k)
frame_vm_group_bin_11484 = frame (4k)
frame_vm_group_bin_11485 = frame (4k)
frame_vm_group_bin_11486 = frame (4k)
frame_vm_group_bin_11487 = frame (4k)
frame_vm_group_bin_11488 = frame (4k)
frame_vm_group_bin_11489 = frame (4k)
frame_vm_group_bin_1149 = frame (4k)
frame_vm_group_bin_11490 = frame (4k)
frame_vm_group_bin_11491 = frame (4k)
frame_vm_group_bin_11492 = frame (4k)
frame_vm_group_bin_11493 = frame (4k)
frame_vm_group_bin_11494 = frame (4k)
frame_vm_group_bin_11495 = frame (4k)
frame_vm_group_bin_11496 = frame (4k)
frame_vm_group_bin_11497 = frame (4k)
frame_vm_group_bin_11498 = frame (4k)
frame_vm_group_bin_11499 = frame (4k)
frame_vm_group_bin_1150 = frame (4k)
frame_vm_group_bin_11500 = frame (4k)
frame_vm_group_bin_11501 = frame (4k)
frame_vm_group_bin_11502 = frame (4k)
frame_vm_group_bin_11503 = frame (4k)
frame_vm_group_bin_11504 = frame (4k)
frame_vm_group_bin_11505 = frame (4k)
frame_vm_group_bin_11506 = frame (4k)
frame_vm_group_bin_11507 = frame (4k)
frame_vm_group_bin_11508 = frame (4k)
frame_vm_group_bin_11509 = frame (4k)
frame_vm_group_bin_1151 = frame (4k)
frame_vm_group_bin_11510 = frame (4k)
frame_vm_group_bin_11511 = frame (4k)
frame_vm_group_bin_11512 = frame (4k)
frame_vm_group_bin_11513 = frame (4k)
frame_vm_group_bin_11514 = frame (4k)
frame_vm_group_bin_11515 = frame (4k)
frame_vm_group_bin_11516 = frame (4k)
frame_vm_group_bin_11517 = frame (4k)
frame_vm_group_bin_11518 = frame (4k)
frame_vm_group_bin_11519 = frame (4k)
frame_vm_group_bin_1152 = frame (4k)
frame_vm_group_bin_11520 = frame (4k)
frame_vm_group_bin_11521 = frame (4k)
frame_vm_group_bin_11522 = frame (4k)
frame_vm_group_bin_11523 = frame (4k)
frame_vm_group_bin_11524 = frame (4k)
frame_vm_group_bin_11525 = frame (4k)
frame_vm_group_bin_11526 = frame (4k)
frame_vm_group_bin_11527 = frame (4k)
frame_vm_group_bin_11528 = frame (4k)
frame_vm_group_bin_11529 = frame (4k)
frame_vm_group_bin_1153 = frame (4k)
frame_vm_group_bin_11530 = frame (4k)
frame_vm_group_bin_11531 = frame (4k)
frame_vm_group_bin_11532 = frame (4k)
frame_vm_group_bin_11533 = frame (4k)
frame_vm_group_bin_11534 = frame (4k)
frame_vm_group_bin_11535 = frame (4k)
frame_vm_group_bin_11536 = frame (4k)
frame_vm_group_bin_11537 = frame (4k)
frame_vm_group_bin_11538 = frame (4k)
frame_vm_group_bin_11539 = frame (4k)
frame_vm_group_bin_1154 = frame (4k)
frame_vm_group_bin_11540 = frame (4k)
frame_vm_group_bin_11541 = frame (4k)
frame_vm_group_bin_11542 = frame (4k)
frame_vm_group_bin_11543 = frame (4k)
frame_vm_group_bin_11544 = frame (4k)
frame_vm_group_bin_11545 = frame (4k)
frame_vm_group_bin_11546 = frame (4k)
frame_vm_group_bin_11547 = frame (4k)
frame_vm_group_bin_11548 = frame (4k)
frame_vm_group_bin_11549 = frame (4k)
frame_vm_group_bin_1155 = frame (4k)
frame_vm_group_bin_11550 = frame (4k)
frame_vm_group_bin_11551 = frame (4k)
frame_vm_group_bin_11552 = frame (4k)
frame_vm_group_bin_11553 = frame (4k)
frame_vm_group_bin_11554 = frame (4k)
frame_vm_group_bin_11555 = frame (4k)
frame_vm_group_bin_11556 = frame (4k)
frame_vm_group_bin_11557 = frame (4k)
frame_vm_group_bin_11558 = frame (4k)
frame_vm_group_bin_11559 = frame (4k)
frame_vm_group_bin_1156 = frame (4k)
frame_vm_group_bin_11560 = frame (4k)
frame_vm_group_bin_11561 = frame (4k)
frame_vm_group_bin_11562 = frame (4k)
frame_vm_group_bin_11563 = frame (4k)
frame_vm_group_bin_11564 = frame (4k)
frame_vm_group_bin_11565 = frame (4k)
frame_vm_group_bin_11566 = frame (4k)
frame_vm_group_bin_11567 = frame (4k)
frame_vm_group_bin_11568 = frame (4k)
frame_vm_group_bin_11569 = frame (4k)
frame_vm_group_bin_1157 = frame (4k)
frame_vm_group_bin_11570 = frame (4k)
frame_vm_group_bin_11571 = frame (4k)
frame_vm_group_bin_11572 = frame (4k)
frame_vm_group_bin_11573 = frame (4k)
frame_vm_group_bin_11574 = frame (4k)
frame_vm_group_bin_11575 = frame (4k)
frame_vm_group_bin_11576 = frame (4k)
frame_vm_group_bin_11577 = frame (4k)
frame_vm_group_bin_11578 = frame (4k)
frame_vm_group_bin_11579 = frame (4k)
frame_vm_group_bin_1158 = frame (4k)
frame_vm_group_bin_11580 = frame (4k)
frame_vm_group_bin_11581 = frame (4k)
frame_vm_group_bin_11582 = frame (4k)
frame_vm_group_bin_11583 = frame (4k)
frame_vm_group_bin_11584 = frame (4k)
frame_vm_group_bin_11585 = frame (4k)
frame_vm_group_bin_11586 = frame (4k)
frame_vm_group_bin_11587 = frame (4k)
frame_vm_group_bin_11588 = frame (4k)
frame_vm_group_bin_11589 = frame (4k)
frame_vm_group_bin_1159 = frame (4k)
frame_vm_group_bin_11590 = frame (4k)
frame_vm_group_bin_11591 = frame (4k)
frame_vm_group_bin_11592 = frame (4k)
frame_vm_group_bin_11593 = frame (4k)
frame_vm_group_bin_11594 = frame (4k)
frame_vm_group_bin_11595 = frame (4k)
frame_vm_group_bin_11596 = frame (4k)
frame_vm_group_bin_11597 = frame (4k)
frame_vm_group_bin_11598 = frame (4k)
frame_vm_group_bin_11599 = frame (4k)
frame_vm_group_bin_1160 = frame (4k)
frame_vm_group_bin_11600 = frame (4k)
frame_vm_group_bin_11601 = frame (4k)
frame_vm_group_bin_11602 = frame (4k)
frame_vm_group_bin_11603 = frame (4k)
frame_vm_group_bin_11604 = frame (4k)
frame_vm_group_bin_11605 = frame (4k)
frame_vm_group_bin_11606 = frame (4k)
frame_vm_group_bin_11607 = frame (4k)
frame_vm_group_bin_11608 = frame (4k)
frame_vm_group_bin_11609 = frame (4k)
frame_vm_group_bin_1161 = frame (4k)
frame_vm_group_bin_11610 = frame (4k)
frame_vm_group_bin_11611 = frame (4k)
frame_vm_group_bin_11612 = frame (4k)
frame_vm_group_bin_11613 = frame (4k)
frame_vm_group_bin_11614 = frame (4k)
frame_vm_group_bin_11615 = frame (4k)
frame_vm_group_bin_11616 = frame (4k)
frame_vm_group_bin_11617 = frame (4k)
frame_vm_group_bin_11618 = frame (4k)
frame_vm_group_bin_11619 = frame (4k)
frame_vm_group_bin_1162 = frame (4k)
frame_vm_group_bin_11620 = frame (4k)
frame_vm_group_bin_11621 = frame (4k)
frame_vm_group_bin_11622 = frame (4k)
frame_vm_group_bin_11623 = frame (4k)
frame_vm_group_bin_11624 = frame (4k)
frame_vm_group_bin_11625 = frame (4k)
frame_vm_group_bin_11626 = frame (4k)
frame_vm_group_bin_11627 = frame (4k)
frame_vm_group_bin_11628 = frame (4k)
frame_vm_group_bin_11629 = frame (4k)
frame_vm_group_bin_1163 = frame (4k)
frame_vm_group_bin_11630 = frame (4k)
frame_vm_group_bin_11631 = frame (4k)
frame_vm_group_bin_11632 = frame (4k)
frame_vm_group_bin_11633 = frame (4k)
frame_vm_group_bin_11634 = frame (4k)
frame_vm_group_bin_11635 = frame (4k)
frame_vm_group_bin_11636 = frame (4k)
frame_vm_group_bin_11637 = frame (4k)
frame_vm_group_bin_11638 = frame (4k)
frame_vm_group_bin_11639 = frame (4k)
frame_vm_group_bin_1164 = frame (4k)
frame_vm_group_bin_11640 = frame (4k)
frame_vm_group_bin_11641 = frame (4k)
frame_vm_group_bin_11642 = frame (4k)
frame_vm_group_bin_11643 = frame (4k)
frame_vm_group_bin_11644 = frame (4k)
frame_vm_group_bin_11645 = frame (4k)
frame_vm_group_bin_11646 = frame (4k)
frame_vm_group_bin_11647 = frame (4k)
frame_vm_group_bin_11648 = frame (4k)
frame_vm_group_bin_11649 = frame (4k)
frame_vm_group_bin_1165 = frame (4k)
frame_vm_group_bin_11650 = frame (4k)
frame_vm_group_bin_11651 = frame (4k)
frame_vm_group_bin_11652 = frame (4k)
frame_vm_group_bin_11653 = frame (4k)
frame_vm_group_bin_11654 = frame (4k)
frame_vm_group_bin_11655 = frame (4k)
frame_vm_group_bin_11656 = frame (4k)
frame_vm_group_bin_11657 = frame (4k)
frame_vm_group_bin_11658 = frame (4k)
frame_vm_group_bin_11659 = frame (4k)
frame_vm_group_bin_1166 = frame (4k)
frame_vm_group_bin_11660 = frame (4k)
frame_vm_group_bin_11661 = frame (4k)
frame_vm_group_bin_11662 = frame (4k)
frame_vm_group_bin_11663 = frame (4k)
frame_vm_group_bin_11664 = frame (4k)
frame_vm_group_bin_11665 = frame (4k)
frame_vm_group_bin_11666 = frame (4k)
frame_vm_group_bin_11667 = frame (4k)
frame_vm_group_bin_11668 = frame (4k)
frame_vm_group_bin_11669 = frame (4k)
frame_vm_group_bin_1167 = frame (4k)
frame_vm_group_bin_11670 = frame (4k)
frame_vm_group_bin_11671 = frame (4k)
frame_vm_group_bin_11672 = frame (4k)
frame_vm_group_bin_11673 = frame (4k)
frame_vm_group_bin_11674 = frame (4k)
frame_vm_group_bin_11675 = frame (4k)
frame_vm_group_bin_11676 = frame (4k)
frame_vm_group_bin_11677 = frame (4k)
frame_vm_group_bin_11678 = frame (4k)
frame_vm_group_bin_11679 = frame (4k)
frame_vm_group_bin_1168 = frame (4k)
frame_vm_group_bin_11680 = frame (4k)
frame_vm_group_bin_11681 = frame (4k)
frame_vm_group_bin_11682 = frame (4k)
frame_vm_group_bin_11683 = frame (4k)
frame_vm_group_bin_11684 = frame (4k)
frame_vm_group_bin_11685 = frame (4k)
frame_vm_group_bin_11686 = frame (4k)
frame_vm_group_bin_11687 = frame (4k)
frame_vm_group_bin_11688 = frame (4k)
frame_vm_group_bin_11689 = frame (4k)
frame_vm_group_bin_1169 = frame (4k)
frame_vm_group_bin_11690 = frame (4k)
frame_vm_group_bin_11691 = frame (4k)
frame_vm_group_bin_11692 = frame (4k)
frame_vm_group_bin_11693 = frame (4k)
frame_vm_group_bin_11694 = frame (4k)
frame_vm_group_bin_11695 = frame (4k)
frame_vm_group_bin_11696 = frame (4k)
frame_vm_group_bin_11697 = frame (4k)
frame_vm_group_bin_11698 = frame (4k)
frame_vm_group_bin_11699 = frame (4k)
frame_vm_group_bin_1170 = frame (4k)
frame_vm_group_bin_11700 = frame (4k)
frame_vm_group_bin_11701 = frame (4k)
frame_vm_group_bin_11702 = frame (4k)
frame_vm_group_bin_11703 = frame (4k)
frame_vm_group_bin_11704 = frame (4k)
frame_vm_group_bin_11705 = frame (4k)
frame_vm_group_bin_11706 = frame (4k)
frame_vm_group_bin_11707 = frame (4k)
frame_vm_group_bin_11708 = frame (4k)
frame_vm_group_bin_11709 = frame (4k)
frame_vm_group_bin_1171 = frame (4k)
frame_vm_group_bin_11710 = frame (4k)
frame_vm_group_bin_11711 = frame (4k)
frame_vm_group_bin_11712 = frame (4k)
frame_vm_group_bin_11713 = frame (4k)
frame_vm_group_bin_11714 = frame (4k)
frame_vm_group_bin_11715 = frame (4k)
frame_vm_group_bin_11716 = frame (4k)
frame_vm_group_bin_11717 = frame (4k)
frame_vm_group_bin_11718 = frame (4k)
frame_vm_group_bin_11719 = frame (4k)
frame_vm_group_bin_1172 = frame (4k)
frame_vm_group_bin_11720 = frame (4k)
frame_vm_group_bin_11721 = frame (4k)
frame_vm_group_bin_11722 = frame (4k)
frame_vm_group_bin_11723 = frame (4k)
frame_vm_group_bin_11724 = frame (4k)
frame_vm_group_bin_11725 = frame (4k)
frame_vm_group_bin_11726 = frame (4k)
frame_vm_group_bin_11727 = frame (4k)
frame_vm_group_bin_11728 = frame (4k)
frame_vm_group_bin_11729 = frame (4k)
frame_vm_group_bin_1173 = frame (4k)
frame_vm_group_bin_11730 = frame (4k)
frame_vm_group_bin_11731 = frame (4k)
frame_vm_group_bin_11732 = frame (4k)
frame_vm_group_bin_11733 = frame (4k)
frame_vm_group_bin_11734 = frame (4k)
frame_vm_group_bin_11735 = frame (4k)
frame_vm_group_bin_11736 = frame (4k)
frame_vm_group_bin_11737 = frame (4k)
frame_vm_group_bin_11738 = frame (4k)
frame_vm_group_bin_11739 = frame (4k)
frame_vm_group_bin_1174 = frame (4k)
frame_vm_group_bin_11740 = frame (4k)
frame_vm_group_bin_11741 = frame (4k)
frame_vm_group_bin_11742 = frame (4k)
frame_vm_group_bin_11743 = frame (4k)
frame_vm_group_bin_11744 = frame (4k)
frame_vm_group_bin_11745 = frame (4k)
frame_vm_group_bin_11746 = frame (4k)
frame_vm_group_bin_11747 = frame (4k)
frame_vm_group_bin_11748 = frame (4k)
frame_vm_group_bin_11749 = frame (4k)
frame_vm_group_bin_1175 = frame (4k)
frame_vm_group_bin_11750 = frame (4k)
frame_vm_group_bin_11751 = frame (4k)
frame_vm_group_bin_11752 = frame (4k)
frame_vm_group_bin_11753 = frame (4k)
frame_vm_group_bin_11754 = frame (4k)
frame_vm_group_bin_11755 = frame (4k)
frame_vm_group_bin_11756 = frame (4k)
frame_vm_group_bin_11757 = frame (4k)
frame_vm_group_bin_11758 = frame (4k)
frame_vm_group_bin_11759 = frame (4k)
frame_vm_group_bin_1176 = frame (4k)
frame_vm_group_bin_11760 = frame (4k)
frame_vm_group_bin_11761 = frame (4k)
frame_vm_group_bin_11762 = frame (4k)
frame_vm_group_bin_11763 = frame (4k)
frame_vm_group_bin_11764 = frame (4k)
frame_vm_group_bin_11765 = frame (4k)
frame_vm_group_bin_11766 = frame (4k)
frame_vm_group_bin_11767 = frame (4k)
frame_vm_group_bin_11768 = frame (4k)
frame_vm_group_bin_11769 = frame (4k)
frame_vm_group_bin_1177 = frame (4k)
frame_vm_group_bin_11770 = frame (4k)
frame_vm_group_bin_11771 = frame (4k)
frame_vm_group_bin_11772 = frame (4k)
frame_vm_group_bin_11773 = frame (4k)
frame_vm_group_bin_11774 = frame (4k)
frame_vm_group_bin_11775 = frame (4k)
frame_vm_group_bin_11776 = frame (4k)
frame_vm_group_bin_11777 = frame (4k)
frame_vm_group_bin_11778 = frame (4k)
frame_vm_group_bin_11779 = frame (4k)
frame_vm_group_bin_1178 = frame (4k)
frame_vm_group_bin_11780 = frame (4k)
frame_vm_group_bin_11781 = frame (4k)
frame_vm_group_bin_11782 = frame (4k)
frame_vm_group_bin_11783 = frame (4k)
frame_vm_group_bin_11784 = frame (4k)
frame_vm_group_bin_11785 = frame (4k)
frame_vm_group_bin_11786 = frame (4k)
frame_vm_group_bin_11787 = frame (4k)
frame_vm_group_bin_11788 = frame (4k)
frame_vm_group_bin_11789 = frame (4k)
frame_vm_group_bin_1179 = frame (4k)
frame_vm_group_bin_11790 = frame (4k)
frame_vm_group_bin_11791 = frame (4k)
frame_vm_group_bin_11792 = frame (4k)
frame_vm_group_bin_11793 = frame (4k)
frame_vm_group_bin_11794 = frame (4k)
frame_vm_group_bin_11795 = frame (4k)
frame_vm_group_bin_11796 = frame (4k)
frame_vm_group_bin_11797 = frame (4k)
frame_vm_group_bin_11798 = frame (4k)
frame_vm_group_bin_11799 = frame (4k)
frame_vm_group_bin_1180 = frame (4k)
frame_vm_group_bin_11800 = frame (4k)
frame_vm_group_bin_11801 = frame (4k)
frame_vm_group_bin_11802 = frame (4k)
frame_vm_group_bin_11803 = frame (4k)
frame_vm_group_bin_11804 = frame (4k)
frame_vm_group_bin_11805 = frame (4k)
frame_vm_group_bin_11806 = frame (4k)
frame_vm_group_bin_11807 = frame (4k)
frame_vm_group_bin_11808 = frame (4k)
frame_vm_group_bin_11809 = frame (4k)
frame_vm_group_bin_1181 = frame (4k)
frame_vm_group_bin_11810 = frame (4k)
frame_vm_group_bin_11811 = frame (4k)
frame_vm_group_bin_11812 = frame (4k)
frame_vm_group_bin_11813 = frame (4k)
frame_vm_group_bin_11814 = frame (4k)
frame_vm_group_bin_11815 = frame (4k)
frame_vm_group_bin_11816 = frame (4k)
frame_vm_group_bin_11817 = frame (4k)
frame_vm_group_bin_11818 = frame (4k)
frame_vm_group_bin_11819 = frame (4k)
frame_vm_group_bin_1182 = frame (4k)
frame_vm_group_bin_11820 = frame (4k)
frame_vm_group_bin_11821 = frame (4k)
frame_vm_group_bin_11822 = frame (4k)
frame_vm_group_bin_11823 = frame (4k)
frame_vm_group_bin_11824 = frame (4k)
frame_vm_group_bin_11825 = frame (4k)
frame_vm_group_bin_11826 = frame (4k)
frame_vm_group_bin_11827 = frame (4k)
frame_vm_group_bin_11828 = frame (4k)
frame_vm_group_bin_11829 = frame (4k)
frame_vm_group_bin_1183 = frame (4k)
frame_vm_group_bin_11830 = frame (4k)
frame_vm_group_bin_11831 = frame (4k)
frame_vm_group_bin_11832 = frame (4k)
frame_vm_group_bin_11833 = frame (4k)
frame_vm_group_bin_11834 = frame (4k)
frame_vm_group_bin_11835 = frame (4k)
frame_vm_group_bin_11836 = frame (4k)
frame_vm_group_bin_11837 = frame (4k)
frame_vm_group_bin_11838 = frame (4k)
frame_vm_group_bin_11839 = frame (4k)
frame_vm_group_bin_1184 = frame (4k)
frame_vm_group_bin_11840 = frame (4k)
frame_vm_group_bin_11841 = frame (4k)
frame_vm_group_bin_11842 = frame (4k)
frame_vm_group_bin_11843 = frame (4k)
frame_vm_group_bin_11844 = frame (4k)
frame_vm_group_bin_11845 = frame (4k)
frame_vm_group_bin_11846 = frame (4k)
frame_vm_group_bin_11847 = frame (4k)
frame_vm_group_bin_11848 = frame (4k)
frame_vm_group_bin_11849 = frame (4k)
frame_vm_group_bin_1185 = frame (4k)
frame_vm_group_bin_11850 = frame (4k)
frame_vm_group_bin_11851 = frame (4k)
frame_vm_group_bin_11852 = frame (4k)
frame_vm_group_bin_11853 = frame (4k)
frame_vm_group_bin_11854 = frame (4k)
frame_vm_group_bin_11855 = frame (4k)
frame_vm_group_bin_11856 = frame (4k)
frame_vm_group_bin_11857 = frame (4k)
frame_vm_group_bin_11858 = frame (4k)
frame_vm_group_bin_11859 = frame (4k)
frame_vm_group_bin_1186 = frame (4k)
frame_vm_group_bin_11860 = frame (4k)
frame_vm_group_bin_11861 = frame (4k)
frame_vm_group_bin_11862 = frame (4k)
frame_vm_group_bin_11863 = frame (4k)
frame_vm_group_bin_11864 = frame (4k)
frame_vm_group_bin_11865 = frame (4k)
frame_vm_group_bin_11866 = frame (4k)
frame_vm_group_bin_11867 = frame (4k)
frame_vm_group_bin_11868 = frame (4k)
frame_vm_group_bin_11869 = frame (4k)
frame_vm_group_bin_1187 = frame (4k)
frame_vm_group_bin_11870 = frame (4k)
frame_vm_group_bin_11871 = frame (4k)
frame_vm_group_bin_11872 = frame (4k)
frame_vm_group_bin_11873 = frame (4k)
frame_vm_group_bin_11874 = frame (4k)
frame_vm_group_bin_11875 = frame (4k)
frame_vm_group_bin_11876 = frame (4k)
frame_vm_group_bin_11877 = frame (4k)
frame_vm_group_bin_11878 = frame (4k)
frame_vm_group_bin_11879 = frame (4k)
frame_vm_group_bin_1188 = frame (4k)
frame_vm_group_bin_11880 = frame (4k)
frame_vm_group_bin_11881 = frame (4k)
frame_vm_group_bin_11882 = frame (4k)
frame_vm_group_bin_11883 = frame (4k)
frame_vm_group_bin_11884 = frame (4k)
frame_vm_group_bin_11885 = frame (4k)
frame_vm_group_bin_11886 = frame (4k)
frame_vm_group_bin_11887 = frame (4k)
frame_vm_group_bin_11888 = frame (4k)
frame_vm_group_bin_11889 = frame (4k)
frame_vm_group_bin_1189 = frame (4k)
frame_vm_group_bin_11890 = frame (4k)
frame_vm_group_bin_11891 = frame (4k)
frame_vm_group_bin_11892 = frame (4k)
frame_vm_group_bin_11893 = frame (4k)
frame_vm_group_bin_11894 = frame (4k)
frame_vm_group_bin_11895 = frame (4k)
frame_vm_group_bin_11896 = frame (4k)
frame_vm_group_bin_11897 = frame (4k)
frame_vm_group_bin_11898 = frame (4k)
frame_vm_group_bin_11899 = frame (4k)
frame_vm_group_bin_1190 = frame (4k)
frame_vm_group_bin_11900 = frame (4k)
frame_vm_group_bin_11901 = frame (4k)
frame_vm_group_bin_11902 = frame (4k)
frame_vm_group_bin_11903 = frame (4k)
frame_vm_group_bin_11904 = frame (4k)
frame_vm_group_bin_11905 = frame (4k)
frame_vm_group_bin_11906 = frame (4k)
frame_vm_group_bin_11907 = frame (4k)
frame_vm_group_bin_11908 = frame (4k)
frame_vm_group_bin_11909 = frame (4k)
frame_vm_group_bin_1191 = frame (4k)
frame_vm_group_bin_11910 = frame (4k)
frame_vm_group_bin_11911 = frame (4k)
frame_vm_group_bin_11912 = frame (4k)
frame_vm_group_bin_11913 = frame (4k)
frame_vm_group_bin_11914 = frame (4k)
frame_vm_group_bin_11915 = frame (4k)
frame_vm_group_bin_11916 = frame (4k)
frame_vm_group_bin_11917 = frame (4k)
frame_vm_group_bin_11918 = frame (4k)
frame_vm_group_bin_11919 = frame (4k)
frame_vm_group_bin_1192 = frame (4k)
frame_vm_group_bin_11920 = frame (4k)
frame_vm_group_bin_11921 = frame (4k)
frame_vm_group_bin_11922 = frame (4k)
frame_vm_group_bin_11923 = frame (4k)
frame_vm_group_bin_11924 = frame (4k)
frame_vm_group_bin_11925 = frame (4k)
frame_vm_group_bin_11926 = frame (4k)
frame_vm_group_bin_11927 = frame (4k)
frame_vm_group_bin_11928 = frame (4k)
frame_vm_group_bin_11929 = frame (4k)
frame_vm_group_bin_1193 = frame (4k)
frame_vm_group_bin_11930 = frame (4k)
frame_vm_group_bin_11931 = frame (4k)
frame_vm_group_bin_11932 = frame (4k)
frame_vm_group_bin_11933 = frame (4k)
frame_vm_group_bin_11934 = frame (4k)
frame_vm_group_bin_11935 = frame (4k)
frame_vm_group_bin_11936 = frame (4k)
frame_vm_group_bin_11937 = frame (4k)
frame_vm_group_bin_11938 = frame (4k)
frame_vm_group_bin_11939 = frame (4k)
frame_vm_group_bin_1194 = frame (4k)
frame_vm_group_bin_11940 = frame (4k)
frame_vm_group_bin_11941 = frame (4k)
frame_vm_group_bin_11942 = frame (4k)
frame_vm_group_bin_11943 = frame (4k)
frame_vm_group_bin_11944 = frame (4k)
frame_vm_group_bin_11945 = frame (4k)
frame_vm_group_bin_11946 = frame (4k)
frame_vm_group_bin_11947 = frame (4k)
frame_vm_group_bin_11948 = frame (4k)
frame_vm_group_bin_11949 = frame (4k)
frame_vm_group_bin_1195 = frame (4k)
frame_vm_group_bin_11950 = frame (4k)
frame_vm_group_bin_11951 = frame (4k)
frame_vm_group_bin_11952 = frame (4k)
frame_vm_group_bin_11953 = frame (4k)
frame_vm_group_bin_11954 = frame (4k)
frame_vm_group_bin_11955 = frame (4k)
frame_vm_group_bin_11956 = frame (4k)
frame_vm_group_bin_11957 = frame (4k)
frame_vm_group_bin_11958 = frame (4k)
frame_vm_group_bin_11959 = frame (4k)
frame_vm_group_bin_1196 = frame (4k)
frame_vm_group_bin_11960 = frame (4k)
frame_vm_group_bin_11961 = frame (4k)
frame_vm_group_bin_11962 = frame (4k)
frame_vm_group_bin_11963 = frame (4k)
frame_vm_group_bin_11964 = frame (4k)
frame_vm_group_bin_11965 = frame (4k)
frame_vm_group_bin_11966 = frame (4k)
frame_vm_group_bin_11967 = frame (4k)
frame_vm_group_bin_11968 = frame (4k)
frame_vm_group_bin_11969 = frame (4k)
frame_vm_group_bin_1197 = frame (4k)
frame_vm_group_bin_11970 = frame (4k)
frame_vm_group_bin_11971 = frame (4k)
frame_vm_group_bin_11972 = frame (4k)
frame_vm_group_bin_11973 = frame (4k)
frame_vm_group_bin_11974 = frame (4k)
frame_vm_group_bin_11975 = frame (4k)
frame_vm_group_bin_11976 = frame (4k)
frame_vm_group_bin_11977 = frame (4k)
frame_vm_group_bin_11978 = frame (4k)
frame_vm_group_bin_11979 = frame (4k)
frame_vm_group_bin_1198 = frame (4k)
frame_vm_group_bin_11980 = frame (4k)
frame_vm_group_bin_11981 = frame (4k)
frame_vm_group_bin_11982 = frame (4k)
frame_vm_group_bin_11983 = frame (4k)
frame_vm_group_bin_11984 = frame (4k)
frame_vm_group_bin_11985 = frame (4k)
frame_vm_group_bin_11986 = frame (4k)
frame_vm_group_bin_11987 = frame (4k)
frame_vm_group_bin_11988 = frame (4k)
frame_vm_group_bin_11989 = frame (4k)
frame_vm_group_bin_1199 = frame (4k)
frame_vm_group_bin_11990 = frame (4k)
frame_vm_group_bin_11991 = frame (4k)
frame_vm_group_bin_11992 = frame (4k)
frame_vm_group_bin_11993 = frame (4k)
frame_vm_group_bin_11994 = frame (4k)
frame_vm_group_bin_11995 = frame (4k)
frame_vm_group_bin_11996 = frame (4k)
frame_vm_group_bin_11997 = frame (4k)
frame_vm_group_bin_11998 = frame (4k)
frame_vm_group_bin_11999 = frame (4k)
frame_vm_group_bin_1200 = frame (4k)
frame_vm_group_bin_12000 = frame (4k)
frame_vm_group_bin_12001 = frame (4k)
frame_vm_group_bin_12002 = frame (4k)
frame_vm_group_bin_12003 = frame (4k)
frame_vm_group_bin_12004 = frame (4k)
frame_vm_group_bin_12005 = frame (4k)
frame_vm_group_bin_12006 = frame (4k)
frame_vm_group_bin_12007 = frame (4k)
frame_vm_group_bin_12008 = frame (4k)
frame_vm_group_bin_12009 = frame (4k)
frame_vm_group_bin_1201 = frame (4k)
frame_vm_group_bin_12010 = frame (4k)
frame_vm_group_bin_12011 = frame (4k)
frame_vm_group_bin_12012 = frame (4k)
frame_vm_group_bin_12013 = frame (4k)
frame_vm_group_bin_12014 = frame (4k)
frame_vm_group_bin_12015 = frame (4k)
frame_vm_group_bin_12016 = frame (4k)
frame_vm_group_bin_12017 = frame (4k)
frame_vm_group_bin_12018 = frame (4k)
frame_vm_group_bin_12019 = frame (4k)
frame_vm_group_bin_1202 = frame (4k)
frame_vm_group_bin_12020 = frame (4k)
frame_vm_group_bin_12021 = frame (4k)
frame_vm_group_bin_12022 = frame (4k)
frame_vm_group_bin_12023 = frame (4k)
frame_vm_group_bin_12024 = frame (4k)
frame_vm_group_bin_12025 = frame (4k)
frame_vm_group_bin_12026 = frame (4k)
frame_vm_group_bin_12027 = frame (4k)
frame_vm_group_bin_12028 = frame (4k)
frame_vm_group_bin_12029 = frame (4k)
frame_vm_group_bin_1203 = frame (4k)
frame_vm_group_bin_12030 = frame (4k)
frame_vm_group_bin_12031 = frame (4k)
frame_vm_group_bin_12032 = frame (4k)
frame_vm_group_bin_12033 = frame (4k)
frame_vm_group_bin_12034 = frame (4k)
frame_vm_group_bin_12035 = frame (4k)
frame_vm_group_bin_12036 = frame (4k)
frame_vm_group_bin_12037 = frame (4k)
frame_vm_group_bin_12038 = frame (4k)
frame_vm_group_bin_12039 = frame (4k)
frame_vm_group_bin_1204 = frame (4k)
frame_vm_group_bin_12040 = frame (4k)
frame_vm_group_bin_12041 = frame (4k)
frame_vm_group_bin_12042 = frame (4k)
frame_vm_group_bin_12043 = frame (4k)
frame_vm_group_bin_12044 = frame (4k)
frame_vm_group_bin_12045 = frame (4k)
frame_vm_group_bin_12046 = frame (4k)
frame_vm_group_bin_12047 = frame (4k)
frame_vm_group_bin_12048 = frame (4k)
frame_vm_group_bin_12049 = frame (4k)
frame_vm_group_bin_1205 = frame (4k)
frame_vm_group_bin_12050 = frame (4k)
frame_vm_group_bin_12051 = frame (4k)
frame_vm_group_bin_12052 = frame (4k)
frame_vm_group_bin_12053 = frame (4k)
frame_vm_group_bin_12054 = frame (4k)
frame_vm_group_bin_12055 = frame (4k)
frame_vm_group_bin_12056 = frame (4k)
frame_vm_group_bin_12057 = frame (4k)
frame_vm_group_bin_12058 = frame (4k)
frame_vm_group_bin_12059 = frame (4k)
frame_vm_group_bin_1206 = frame (4k)
frame_vm_group_bin_12060 = frame (4k)
frame_vm_group_bin_12061 = frame (4k)
frame_vm_group_bin_12062 = frame (4k)
frame_vm_group_bin_12063 = frame (4k)
frame_vm_group_bin_12064 = frame (4k)
frame_vm_group_bin_12065 = frame (4k)
frame_vm_group_bin_12066 = frame (4k)
frame_vm_group_bin_12067 = frame (4k)
frame_vm_group_bin_12068 = frame (4k)
frame_vm_group_bin_12069 = frame (4k)
frame_vm_group_bin_1207 = frame (4k)
frame_vm_group_bin_12070 = frame (4k)
frame_vm_group_bin_12071 = frame (4k)
frame_vm_group_bin_12072 = frame (4k)
frame_vm_group_bin_12073 = frame (4k)
frame_vm_group_bin_12074 = frame (4k)
frame_vm_group_bin_12075 = frame (4k)
frame_vm_group_bin_12076 = frame (4k)
frame_vm_group_bin_12077 = frame (4k)
frame_vm_group_bin_12078 = frame (4k)
frame_vm_group_bin_12079 = frame (4k)
frame_vm_group_bin_1208 = frame (4k)
frame_vm_group_bin_12080 = frame (4k)
frame_vm_group_bin_12081 = frame (4k)
frame_vm_group_bin_12082 = frame (4k)
frame_vm_group_bin_12083 = frame (4k)
frame_vm_group_bin_12084 = frame (4k)
frame_vm_group_bin_12085 = frame (4k)
frame_vm_group_bin_12086 = frame (4k)
frame_vm_group_bin_12087 = frame (4k)
frame_vm_group_bin_12088 = frame (4k)
frame_vm_group_bin_12089 = frame (4k)
frame_vm_group_bin_1209 = frame (4k)
frame_vm_group_bin_12090 = frame (4k)
frame_vm_group_bin_12091 = frame (4k)
frame_vm_group_bin_12092 = frame (4k)
frame_vm_group_bin_12093 = frame (4k)
frame_vm_group_bin_12094 = frame (4k)
frame_vm_group_bin_12095 = frame (4k)
frame_vm_group_bin_12096 = frame (4k)
frame_vm_group_bin_12097 = frame (4k)
frame_vm_group_bin_12098 = frame (4k)
frame_vm_group_bin_12099 = frame (4k)
frame_vm_group_bin_1210 = frame (4k)
frame_vm_group_bin_12100 = frame (4k)
frame_vm_group_bin_12101 = frame (4k)
frame_vm_group_bin_12102 = frame (4k)
frame_vm_group_bin_12103 = frame (4k)
frame_vm_group_bin_12104 = frame (4k)
frame_vm_group_bin_12105 = frame (4k)
frame_vm_group_bin_12106 = frame (4k)
frame_vm_group_bin_12107 = frame (4k)
frame_vm_group_bin_12108 = frame (4k)
frame_vm_group_bin_12109 = frame (4k)
frame_vm_group_bin_1211 = frame (4k)
frame_vm_group_bin_12110 = frame (4k)
frame_vm_group_bin_12111 = frame (4k)
frame_vm_group_bin_12112 = frame (4k)
frame_vm_group_bin_12113 = frame (4k)
frame_vm_group_bin_12114 = frame (4k)
frame_vm_group_bin_12115 = frame (4k)
frame_vm_group_bin_12116 = frame (4k)
frame_vm_group_bin_12117 = frame (4k)
frame_vm_group_bin_12118 = frame (4k)
frame_vm_group_bin_12119 = frame (4k)
frame_vm_group_bin_1212 = frame (4k)
frame_vm_group_bin_12120 = frame (4k)
frame_vm_group_bin_12121 = frame (4k)
frame_vm_group_bin_12122 = frame (4k)
frame_vm_group_bin_12123 = frame (4k)
frame_vm_group_bin_12124 = frame (4k)
frame_vm_group_bin_12125 = frame (4k)
frame_vm_group_bin_12126 = frame (4k)
frame_vm_group_bin_12127 = frame (4k)
frame_vm_group_bin_12128 = frame (4k)
frame_vm_group_bin_12129 = frame (4k)
frame_vm_group_bin_1213 = frame (4k)
frame_vm_group_bin_12130 = frame (4k)
frame_vm_group_bin_12131 = frame (4k)
frame_vm_group_bin_12132 = frame (4k)
frame_vm_group_bin_12133 = frame (4k)
frame_vm_group_bin_12134 = frame (4k)
frame_vm_group_bin_12135 = frame (4k)
frame_vm_group_bin_12136 = frame (4k)
frame_vm_group_bin_12137 = frame (4k)
frame_vm_group_bin_12138 = frame (4k)
frame_vm_group_bin_12139 = frame (4k)
frame_vm_group_bin_1214 = frame (4k)
frame_vm_group_bin_12140 = frame (4k)
frame_vm_group_bin_12141 = frame (4k)
frame_vm_group_bin_12142 = frame (4k)
frame_vm_group_bin_12143 = frame (4k)
frame_vm_group_bin_12144 = frame (4k)
frame_vm_group_bin_12145 = frame (4k)
frame_vm_group_bin_12146 = frame (4k)
frame_vm_group_bin_12147 = frame (4k)
frame_vm_group_bin_12148 = frame (4k)
frame_vm_group_bin_12149 = frame (4k)
frame_vm_group_bin_1215 = frame (4k)
frame_vm_group_bin_12150 = frame (4k)
frame_vm_group_bin_12151 = frame (4k)
frame_vm_group_bin_12152 = frame (4k)
frame_vm_group_bin_12153 = frame (4k)
frame_vm_group_bin_12154 = frame (4k)
frame_vm_group_bin_12155 = frame (4k)
frame_vm_group_bin_12156 = frame (4k)
frame_vm_group_bin_12157 = frame (4k)
frame_vm_group_bin_12158 = frame (4k)
frame_vm_group_bin_12159 = frame (4k)
frame_vm_group_bin_1216 = frame (4k)
frame_vm_group_bin_12160 = frame (4k)
frame_vm_group_bin_12161 = frame (4k)
frame_vm_group_bin_12162 = frame (4k)
frame_vm_group_bin_12163 = frame (4k)
frame_vm_group_bin_12164 = frame (4k)
frame_vm_group_bin_12165 = frame (4k)
frame_vm_group_bin_12166 = frame (4k)
frame_vm_group_bin_12167 = frame (4k)
frame_vm_group_bin_12168 = frame (4k)
frame_vm_group_bin_12169 = frame (4k)
frame_vm_group_bin_1217 = frame (4k)
frame_vm_group_bin_12170 = frame (4k)
frame_vm_group_bin_12171 = frame (4k)
frame_vm_group_bin_12172 = frame (4k)
frame_vm_group_bin_12173 = frame (4k)
frame_vm_group_bin_12174 = frame (4k)
frame_vm_group_bin_12175 = frame (4k)
frame_vm_group_bin_12176 = frame (4k)
frame_vm_group_bin_12177 = frame (4k)
frame_vm_group_bin_12178 = frame (4k)
frame_vm_group_bin_12179 = frame (4k)
frame_vm_group_bin_1218 = frame (4k)
frame_vm_group_bin_12180 = frame (4k)
frame_vm_group_bin_12181 = frame (4k)
frame_vm_group_bin_12182 = frame (4k)
frame_vm_group_bin_12183 = frame (4k)
frame_vm_group_bin_12184 = frame (4k)
frame_vm_group_bin_12185 = frame (4k)
frame_vm_group_bin_12186 = frame (4k)
frame_vm_group_bin_12187 = frame (4k)
frame_vm_group_bin_12188 = frame (4k)
frame_vm_group_bin_12189 = frame (4k)
frame_vm_group_bin_1219 = frame (4k)
frame_vm_group_bin_12190 = frame (4k)
frame_vm_group_bin_12191 = frame (4k)
frame_vm_group_bin_12192 = frame (4k)
frame_vm_group_bin_12193 = frame (4k)
frame_vm_group_bin_12194 = frame (4k)
frame_vm_group_bin_12195 = frame (4k)
frame_vm_group_bin_12196 = frame (4k)
frame_vm_group_bin_12197 = frame (4k)
frame_vm_group_bin_12198 = frame (4k)
frame_vm_group_bin_12199 = frame (4k)
frame_vm_group_bin_1220 = frame (4k)
frame_vm_group_bin_12200 = frame (4k)
frame_vm_group_bin_12201 = frame (4k)
frame_vm_group_bin_12202 = frame (4k)
frame_vm_group_bin_12203 = frame (4k)
frame_vm_group_bin_12204 = frame (4k)
frame_vm_group_bin_12205 = frame (4k)
frame_vm_group_bin_12206 = frame (4k)
frame_vm_group_bin_12207 = frame (4k)
frame_vm_group_bin_12208 = frame (4k)
frame_vm_group_bin_12209 = frame (4k)
frame_vm_group_bin_1221 = frame (4k)
frame_vm_group_bin_12210 = frame (4k)
frame_vm_group_bin_12211 = frame (4k)
frame_vm_group_bin_12212 = frame (4k)
frame_vm_group_bin_12213 = frame (4k)
frame_vm_group_bin_12214 = frame (4k)
frame_vm_group_bin_12215 = frame (4k)
frame_vm_group_bin_12216 = frame (4k)
frame_vm_group_bin_12217 = frame (4k)
frame_vm_group_bin_12218 = frame (4k)
frame_vm_group_bin_12219 = frame (4k)
frame_vm_group_bin_1222 = frame (4k)
frame_vm_group_bin_12220 = frame (4k)
frame_vm_group_bin_12221 = frame (4k)
frame_vm_group_bin_12222 = frame (4k)
frame_vm_group_bin_12223 = frame (4k)
frame_vm_group_bin_12224 = frame (4k)
frame_vm_group_bin_12225 = frame (4k)
frame_vm_group_bin_12226 = frame (4k)
frame_vm_group_bin_12227 = frame (4k)
frame_vm_group_bin_12228 = frame (4k)
frame_vm_group_bin_12229 = frame (4k)
frame_vm_group_bin_1223 = frame (4k)
frame_vm_group_bin_12230 = frame (4k)
frame_vm_group_bin_12231 = frame (4k)
frame_vm_group_bin_12232 = frame (4k)
frame_vm_group_bin_12233 = frame (4k)
frame_vm_group_bin_12234 = frame (4k)
frame_vm_group_bin_12235 = frame (4k)
frame_vm_group_bin_12236 = frame (4k)
frame_vm_group_bin_12237 = frame (4k)
frame_vm_group_bin_12238 = frame (4k)
frame_vm_group_bin_12239 = frame (4k)
frame_vm_group_bin_1224 = frame (4k)
frame_vm_group_bin_12240 = frame (4k)
frame_vm_group_bin_12241 = frame (4k)
frame_vm_group_bin_12242 = frame (4k)
frame_vm_group_bin_12243 = frame (4k)
frame_vm_group_bin_12244 = frame (4k)
frame_vm_group_bin_12245 = frame (4k)
frame_vm_group_bin_12246 = frame (4k)
frame_vm_group_bin_12247 = frame (4k)
frame_vm_group_bin_12248 = frame (4k)
frame_vm_group_bin_12249 = frame (4k)
frame_vm_group_bin_1225 = frame (4k)
frame_vm_group_bin_12250 = frame (4k)
frame_vm_group_bin_12251 = frame (4k)
frame_vm_group_bin_12252 = frame (4k)
frame_vm_group_bin_12253 = frame (4k)
frame_vm_group_bin_12254 = frame (4k)
frame_vm_group_bin_12255 = frame (4k)
frame_vm_group_bin_12256 = frame (4k)
frame_vm_group_bin_12257 = frame (4k)
frame_vm_group_bin_12258 = frame (4k)
frame_vm_group_bin_12259 = frame (4k)
frame_vm_group_bin_1226 = frame (4k)
frame_vm_group_bin_12260 = frame (4k)
frame_vm_group_bin_12261 = frame (4k)
frame_vm_group_bin_12262 = frame (4k)
frame_vm_group_bin_12263 = frame (4k)
frame_vm_group_bin_12264 = frame (4k)
frame_vm_group_bin_12265 = frame (4k)
frame_vm_group_bin_12266 = frame (4k)
frame_vm_group_bin_12267 = frame (4k)
frame_vm_group_bin_12268 = frame (4k)
frame_vm_group_bin_12269 = frame (4k)
frame_vm_group_bin_1227 = frame (4k)
frame_vm_group_bin_12270 = frame (4k)
frame_vm_group_bin_12271 = frame (4k)
frame_vm_group_bin_12272 = frame (4k)
frame_vm_group_bin_12273 = frame (4k)
frame_vm_group_bin_12274 = frame (4k)
frame_vm_group_bin_12275 = frame (4k)
frame_vm_group_bin_12276 = frame (4k)
frame_vm_group_bin_12277 = frame (4k)
frame_vm_group_bin_12278 = frame (4k)
frame_vm_group_bin_12279 = frame (4k)
frame_vm_group_bin_1228 = frame (4k)
frame_vm_group_bin_12280 = frame (4k)
frame_vm_group_bin_12281 = frame (4k)
frame_vm_group_bin_12282 = frame (4k)
frame_vm_group_bin_12283 = frame (4k)
frame_vm_group_bin_12284 = frame (4k)
frame_vm_group_bin_12285 = frame (4k)
frame_vm_group_bin_12286 = frame (4k)
frame_vm_group_bin_12287 = frame (4k)
frame_vm_group_bin_12288 = frame (4k)
frame_vm_group_bin_12289 = frame (4k)
frame_vm_group_bin_1229 = frame (4k)
frame_vm_group_bin_12290 = frame (4k)
frame_vm_group_bin_12291 = frame (4k)
frame_vm_group_bin_12292 = frame (4k)
frame_vm_group_bin_12293 = frame (4k)
frame_vm_group_bin_12294 = frame (4k)
frame_vm_group_bin_12295 = frame (4k)
frame_vm_group_bin_12296 = frame (4k)
frame_vm_group_bin_12297 = frame (4k)
frame_vm_group_bin_12298 = frame (4k)
frame_vm_group_bin_12299 = frame (4k)
frame_vm_group_bin_1230 = frame (4k)
frame_vm_group_bin_12300 = frame (4k)
frame_vm_group_bin_12301 = frame (4k)
frame_vm_group_bin_12302 = frame (4k)
frame_vm_group_bin_12303 = frame (4k)
frame_vm_group_bin_12304 = frame (4k)
frame_vm_group_bin_12305 = frame (4k)
frame_vm_group_bin_12306 = frame (4k)
frame_vm_group_bin_12307 = frame (4k)
frame_vm_group_bin_12308 = frame (4k)
frame_vm_group_bin_12309 = frame (4k)
frame_vm_group_bin_1231 = frame (4k)
frame_vm_group_bin_12310 = frame (4k)
frame_vm_group_bin_12311 = frame (4k)
frame_vm_group_bin_12312 = frame (4k)
frame_vm_group_bin_12313 = frame (4k)
frame_vm_group_bin_12314 = frame (4k)
frame_vm_group_bin_12315 = frame (4k)
frame_vm_group_bin_12316 = frame (4k)
frame_vm_group_bin_12317 = frame (4k)
frame_vm_group_bin_12318 = frame (4k)
frame_vm_group_bin_12319 = frame (4k)
frame_vm_group_bin_1232 = frame (4k)
frame_vm_group_bin_12320 = frame (4k)
frame_vm_group_bin_12321 = frame (4k)
frame_vm_group_bin_12322 = frame (4k)
frame_vm_group_bin_12323 = frame (4k)
frame_vm_group_bin_12324 = frame (4k)
frame_vm_group_bin_12325 = frame (4k)
frame_vm_group_bin_12326 = frame (4k)
frame_vm_group_bin_12327 = frame (4k)
frame_vm_group_bin_12328 = frame (4k)
frame_vm_group_bin_12329 = frame (4k)
frame_vm_group_bin_1233 = frame (4k)
frame_vm_group_bin_12330 = frame (4k)
frame_vm_group_bin_12331 = frame (4k)
frame_vm_group_bin_12332 = frame (4k)
frame_vm_group_bin_12333 = frame (4k)
frame_vm_group_bin_12334 = frame (4k)
frame_vm_group_bin_12335 = frame (4k)
frame_vm_group_bin_12336 = frame (4k)
frame_vm_group_bin_12337 = frame (4k)
frame_vm_group_bin_12338 = frame (4k)
frame_vm_group_bin_12339 = frame (4k)
frame_vm_group_bin_1234 = frame (4k)
frame_vm_group_bin_12340 = frame (4k)
frame_vm_group_bin_12341 = frame (4k)
frame_vm_group_bin_12342 = frame (4k)
frame_vm_group_bin_12343 = frame (4k)
frame_vm_group_bin_12344 = frame (4k)
frame_vm_group_bin_12345 = frame (4k)
frame_vm_group_bin_12346 = frame (4k)
frame_vm_group_bin_12347 = frame (4k)
frame_vm_group_bin_12348 = frame (4k)
frame_vm_group_bin_12349 = frame (4k)
frame_vm_group_bin_1235 = frame (4k)
frame_vm_group_bin_12350 = frame (4k)
frame_vm_group_bin_12352 = frame (4k)
frame_vm_group_bin_12353 = frame (4k)
frame_vm_group_bin_12354 = frame (4k)
frame_vm_group_bin_12355 = frame (4k)
frame_vm_group_bin_12356 = frame (4k)
frame_vm_group_bin_12357 = frame (4k)
frame_vm_group_bin_12358 = frame (4k)
frame_vm_group_bin_12359 = frame (4k)
frame_vm_group_bin_1236 = frame (4k)
frame_vm_group_bin_12360 = frame (4k)
frame_vm_group_bin_12361 = frame (4k)
frame_vm_group_bin_12362 = frame (4k)
frame_vm_group_bin_12363 = frame (4k)
frame_vm_group_bin_12364 = frame (4k)
frame_vm_group_bin_12365 = frame (4k)
frame_vm_group_bin_12366 = frame (4k)
frame_vm_group_bin_12367 = frame (4k)
frame_vm_group_bin_12368 = frame (4k)
frame_vm_group_bin_12369 = frame (4k)
frame_vm_group_bin_1237 = frame (4k)
frame_vm_group_bin_12370 = frame (4k)
frame_vm_group_bin_12371 = frame (4k)
frame_vm_group_bin_12372 = frame (4k)
frame_vm_group_bin_12373 = frame (4k)
frame_vm_group_bin_12374 = frame (4k)
frame_vm_group_bin_12375 = frame (4k)
frame_vm_group_bin_12376 = frame (4k)
frame_vm_group_bin_12377 = frame (4k)
frame_vm_group_bin_12378 = frame (4k)
frame_vm_group_bin_12379 = frame (4k)
frame_vm_group_bin_1238 = frame (4k)
frame_vm_group_bin_12380 = frame (4k)
frame_vm_group_bin_12381 = frame (4k)
frame_vm_group_bin_12382 = frame (4k)
frame_vm_group_bin_12383 = frame (4k)
frame_vm_group_bin_12384 = frame (4k)
frame_vm_group_bin_12385 = frame (4k)
frame_vm_group_bin_12386 = frame (4k)
frame_vm_group_bin_12387 = frame (4k)
frame_vm_group_bin_12388 = frame (4k)
frame_vm_group_bin_12389 = frame (4k)
frame_vm_group_bin_1239 = frame (4k)
frame_vm_group_bin_12390 = frame (4k)
frame_vm_group_bin_12391 = frame (4k)
frame_vm_group_bin_12392 = frame (4k)
frame_vm_group_bin_12393 = frame (4k)
frame_vm_group_bin_12394 = frame (4k)
frame_vm_group_bin_12395 = frame (4k)
frame_vm_group_bin_12396 = frame (4k)
frame_vm_group_bin_12397 = frame (4k)
frame_vm_group_bin_12398 = frame (4k)
frame_vm_group_bin_12399 = frame (4k)
frame_vm_group_bin_1240 = frame (4k)
frame_vm_group_bin_12400 = frame (4k)
frame_vm_group_bin_12401 = frame (4k)
frame_vm_group_bin_12402 = frame (4k)
frame_vm_group_bin_12403 = frame (4k)
frame_vm_group_bin_12404 = frame (4k)
frame_vm_group_bin_12405 = frame (4k)
frame_vm_group_bin_12406 = frame (4k)
frame_vm_group_bin_12407 = frame (4k)
frame_vm_group_bin_12408 = frame (4k)
frame_vm_group_bin_12409 = frame (4k)
frame_vm_group_bin_1241 = frame (4k)
frame_vm_group_bin_12410 = frame (4k)
frame_vm_group_bin_12411 = frame (4k)
frame_vm_group_bin_12412 = frame (4k)
frame_vm_group_bin_12413 = frame (4k)
frame_vm_group_bin_12414 = frame (4k)
frame_vm_group_bin_12415 = frame (4k)
frame_vm_group_bin_12416 = frame (4k)
frame_vm_group_bin_12418 = frame (4k)
frame_vm_group_bin_12419 = frame (4k)
frame_vm_group_bin_1242 = frame (4k)
frame_vm_group_bin_12420 = frame (4k)
frame_vm_group_bin_12421 = frame (4k)
frame_vm_group_bin_12422 = frame (4k)
frame_vm_group_bin_12423 = frame (4k)
frame_vm_group_bin_12424 = frame (4k)
frame_vm_group_bin_12425 = frame (4k)
frame_vm_group_bin_12426 = frame (4k)
frame_vm_group_bin_12427 = frame (4k)
frame_vm_group_bin_12428 = frame (4k)
frame_vm_group_bin_12429 = frame (4k)
frame_vm_group_bin_1243 = frame (4k)
frame_vm_group_bin_12430 = frame (4k)
frame_vm_group_bin_12431 = frame (4k)
frame_vm_group_bin_12432 = frame (4k)
frame_vm_group_bin_12433 = frame (4k)
frame_vm_group_bin_12434 = frame (4k)
frame_vm_group_bin_12435 = frame (4k)
frame_vm_group_bin_12436 = frame (4k)
frame_vm_group_bin_12437 = frame (4k)
frame_vm_group_bin_12438 = frame (4k)
frame_vm_group_bin_12439 = frame (4k)
frame_vm_group_bin_1244 = frame (4k)
frame_vm_group_bin_12440 = frame (4k)
frame_vm_group_bin_12441 = frame (4k)
frame_vm_group_bin_12442 = frame (4k)
frame_vm_group_bin_12443 = frame (4k)
frame_vm_group_bin_12444 = frame (4k)
frame_vm_group_bin_12445 = frame (4k)
frame_vm_group_bin_12446 = frame (4k)
frame_vm_group_bin_12447 = frame (4k)
frame_vm_group_bin_12448 = frame (4k)
frame_vm_group_bin_12449 = frame (4k)
frame_vm_group_bin_1245 = frame (4k)
frame_vm_group_bin_12450 = frame (4k)
frame_vm_group_bin_12451 = frame (4k)
frame_vm_group_bin_12452 = frame (4k)
frame_vm_group_bin_12453 = frame (4k)
frame_vm_group_bin_12454 = frame (4k)
frame_vm_group_bin_12455 = frame (4k)
frame_vm_group_bin_12456 = frame (4k)
frame_vm_group_bin_12457 = frame (4k)
frame_vm_group_bin_12458 = frame (4k)
frame_vm_group_bin_12459 = frame (4k)
frame_vm_group_bin_1246 = frame (4k)
frame_vm_group_bin_12460 = frame (4k)
frame_vm_group_bin_12461 = frame (4k)
frame_vm_group_bin_12462 = frame (4k)
frame_vm_group_bin_12463 = frame (4k)
frame_vm_group_bin_12464 = frame (4k)
frame_vm_group_bin_12465 = frame (4k)
frame_vm_group_bin_12466 = frame (4k)
frame_vm_group_bin_12467 = frame (4k)
frame_vm_group_bin_12468 = frame (4k)
frame_vm_group_bin_12469 = frame (4k)
frame_vm_group_bin_1247 = frame (4k)
frame_vm_group_bin_12470 = frame (4k)
frame_vm_group_bin_12471 = frame (4k)
frame_vm_group_bin_12472 = frame (4k)
frame_vm_group_bin_12473 = frame (4k)
frame_vm_group_bin_12474 = frame (4k)
frame_vm_group_bin_12475 = frame (4k)
frame_vm_group_bin_12476 = frame (4k)
frame_vm_group_bin_12477 = frame (4k)
frame_vm_group_bin_12478 = frame (4k)
frame_vm_group_bin_12479 = frame (4k)
frame_vm_group_bin_1248 = frame (4k)
frame_vm_group_bin_12480 = frame (4k)
frame_vm_group_bin_12481 = frame (4k)
frame_vm_group_bin_12482 = frame (4k)
frame_vm_group_bin_12483 = frame (4k)
frame_vm_group_bin_12484 = frame (4k)
frame_vm_group_bin_12485 = frame (4k)
frame_vm_group_bin_12486 = frame (4k)
frame_vm_group_bin_12487 = frame (4k)
frame_vm_group_bin_12488 = frame (4k)
frame_vm_group_bin_12489 = frame (4k)
frame_vm_group_bin_1249 = frame (4k)
frame_vm_group_bin_12490 = frame (4k)
frame_vm_group_bin_12491 = frame (4k)
frame_vm_group_bin_12492 = frame (4k)
frame_vm_group_bin_12493 = frame (4k)
frame_vm_group_bin_12494 = frame (4k)
frame_vm_group_bin_12495 = frame (4k)
frame_vm_group_bin_12496 = frame (4k)
frame_vm_group_bin_12497 = frame (4k)
frame_vm_group_bin_12498 = frame (4k)
frame_vm_group_bin_12499 = frame (4k)
frame_vm_group_bin_1250 = frame (4k)
frame_vm_group_bin_12500 = frame (4k)
frame_vm_group_bin_12501 = frame (4k)
frame_vm_group_bin_12502 = frame (4k)
frame_vm_group_bin_12503 = frame (4k)
frame_vm_group_bin_12504 = frame (4k)
frame_vm_group_bin_12505 = frame (4k)
frame_vm_group_bin_12506 = frame (4k)
frame_vm_group_bin_12507 = frame (4k)
frame_vm_group_bin_12508 = frame (4k)
frame_vm_group_bin_12509 = frame (4k)
frame_vm_group_bin_1251 = frame (4k)
frame_vm_group_bin_12510 = frame (4k)
frame_vm_group_bin_12511 = frame (4k)
frame_vm_group_bin_12512 = frame (4k)
frame_vm_group_bin_12513 = frame (4k)
frame_vm_group_bin_12514 = frame (4k)
frame_vm_group_bin_12515 = frame (4k)
frame_vm_group_bin_12516 = frame (4k)
frame_vm_group_bin_12517 = frame (4k)
frame_vm_group_bin_12518 = frame (4k)
frame_vm_group_bin_12519 = frame (4k)
frame_vm_group_bin_1252 = frame (4k)
frame_vm_group_bin_12520 = frame (4k)
frame_vm_group_bin_12521 = frame (4k)
frame_vm_group_bin_12522 = frame (4k)
frame_vm_group_bin_12523 = frame (4k)
frame_vm_group_bin_12524 = frame (4k)
frame_vm_group_bin_12525 = frame (4k)
frame_vm_group_bin_12526 = frame (4k)
frame_vm_group_bin_12527 = frame (4k)
frame_vm_group_bin_12528 = frame (4k)
frame_vm_group_bin_12529 = frame (4k)
frame_vm_group_bin_1253 = frame (4k)
frame_vm_group_bin_12530 = frame (4k)
frame_vm_group_bin_12531 = frame (4k)
frame_vm_group_bin_12532 = frame (4k)
frame_vm_group_bin_12533 = frame (4k)
frame_vm_group_bin_12534 = frame (4k)
frame_vm_group_bin_12535 = frame (4k)
frame_vm_group_bin_12536 = frame (4k)
frame_vm_group_bin_12537 = frame (4k)
frame_vm_group_bin_12538 = frame (4k)
frame_vm_group_bin_12539 = frame (4k)
frame_vm_group_bin_1254 = frame (4k)
frame_vm_group_bin_12540 = frame (4k)
frame_vm_group_bin_12541 = frame (4k)
frame_vm_group_bin_12542 = frame (4k)
frame_vm_group_bin_12543 = frame (4k)
frame_vm_group_bin_12544 = frame (4k)
frame_vm_group_bin_12545 = frame (4k)
frame_vm_group_bin_12546 = frame (4k)
frame_vm_group_bin_12547 = frame (4k)
frame_vm_group_bin_12548 = frame (4k)
frame_vm_group_bin_12549 = frame (4k)
frame_vm_group_bin_1255 = frame (4k)
frame_vm_group_bin_12550 = frame (4k)
frame_vm_group_bin_12551 = frame (4k)
frame_vm_group_bin_12552 = frame (4k)
frame_vm_group_bin_12553 = frame (4k)
frame_vm_group_bin_12554 = frame (4k)
frame_vm_group_bin_12555 = frame (4k)
frame_vm_group_bin_12556 = frame (4k)
frame_vm_group_bin_12557 = frame (4k)
frame_vm_group_bin_12558 = frame (4k)
frame_vm_group_bin_12559 = frame (4k)
frame_vm_group_bin_1256 = frame (4k)
frame_vm_group_bin_12560 = frame (4k)
frame_vm_group_bin_12561 = frame (4k)
frame_vm_group_bin_12562 = frame (4k)
frame_vm_group_bin_12563 = frame (4k)
frame_vm_group_bin_12564 = frame (4k)
frame_vm_group_bin_12565 = frame (4k)
frame_vm_group_bin_12566 = frame (4k)
frame_vm_group_bin_12567 = frame (4k)
frame_vm_group_bin_12568 = frame (4k)
frame_vm_group_bin_12569 = frame (4k)
frame_vm_group_bin_1257 = frame (4k)
frame_vm_group_bin_12570 = frame (4k)
frame_vm_group_bin_12571 = frame (4k)
frame_vm_group_bin_12572 = frame (4k)
frame_vm_group_bin_12573 = frame (4k)
frame_vm_group_bin_12574 = frame (4k)
frame_vm_group_bin_12575 = frame (4k)
frame_vm_group_bin_12576 = frame (4k)
frame_vm_group_bin_12577 = frame (4k)
frame_vm_group_bin_12578 = frame (4k)
frame_vm_group_bin_12579 = frame (4k)
frame_vm_group_bin_1258 = frame (4k)
frame_vm_group_bin_12580 = frame (4k)
frame_vm_group_bin_12581 = frame (4k)
frame_vm_group_bin_12582 = frame (4k)
frame_vm_group_bin_12583 = frame (4k)
frame_vm_group_bin_12584 = frame (4k)
frame_vm_group_bin_12585 = frame (4k)
frame_vm_group_bin_12586 = frame (4k)
frame_vm_group_bin_12587 = frame (4k)
frame_vm_group_bin_12588 = frame (4k)
frame_vm_group_bin_12589 = frame (4k)
frame_vm_group_bin_1259 = frame (4k)
frame_vm_group_bin_12590 = frame (4k)
frame_vm_group_bin_12591 = frame (4k)
frame_vm_group_bin_12592 = frame (4k)
frame_vm_group_bin_12593 = frame (4k)
frame_vm_group_bin_12594 = frame (4k)
frame_vm_group_bin_12595 = frame (4k)
frame_vm_group_bin_12596 = frame (4k)
frame_vm_group_bin_12597 = frame (4k)
frame_vm_group_bin_12598 = frame (4k)
frame_vm_group_bin_12599 = frame (4k)
frame_vm_group_bin_1260 = frame (4k)
frame_vm_group_bin_12600 = frame (4k)
frame_vm_group_bin_12601 = frame (4k)
frame_vm_group_bin_12602 = frame (4k)
frame_vm_group_bin_12603 = frame (4k)
frame_vm_group_bin_12604 = frame (4k)
frame_vm_group_bin_12605 = frame (4k)
frame_vm_group_bin_12606 = frame (4k)
frame_vm_group_bin_12607 = frame (4k)
frame_vm_group_bin_12608 = frame (4k)
frame_vm_group_bin_12609 = frame (4k)
frame_vm_group_bin_1261 = frame (4k)
frame_vm_group_bin_12610 = frame (4k)
frame_vm_group_bin_12611 = frame (4k)
frame_vm_group_bin_12612 = frame (4k)
frame_vm_group_bin_12613 = frame (4k)
frame_vm_group_bin_12614 = frame (4k)
frame_vm_group_bin_12615 = frame (4k)
frame_vm_group_bin_12616 = frame (4k)
frame_vm_group_bin_12617 = frame (4k)
frame_vm_group_bin_12618 = frame (4k)
frame_vm_group_bin_12619 = frame (4k)
frame_vm_group_bin_1262 = frame (4k)
frame_vm_group_bin_12620 = frame (4k)
frame_vm_group_bin_12621 = frame (4k)
frame_vm_group_bin_12622 = frame (4k)
frame_vm_group_bin_12623 = frame (4k)
frame_vm_group_bin_12624 = frame (4k)
frame_vm_group_bin_12625 = frame (4k)
frame_vm_group_bin_12626 = frame (4k)
frame_vm_group_bin_12627 = frame (4k)
frame_vm_group_bin_12628 = frame (4k)
frame_vm_group_bin_12629 = frame (4k)
frame_vm_group_bin_1263 = frame (4k)
frame_vm_group_bin_12630 = frame (4k)
frame_vm_group_bin_12631 = frame (4k)
frame_vm_group_bin_12632 = frame (4k)
frame_vm_group_bin_12633 = frame (4k)
frame_vm_group_bin_12634 = frame (4k)
frame_vm_group_bin_12635 = frame (4k)
frame_vm_group_bin_12636 = frame (4k)
frame_vm_group_bin_12637 = frame (4k)
frame_vm_group_bin_12638 = frame (4k)
frame_vm_group_bin_12639 = frame (4k)
frame_vm_group_bin_1264 = frame (4k)
frame_vm_group_bin_12640 = frame (4k)
frame_vm_group_bin_12641 = frame (4k)
frame_vm_group_bin_12642 = frame (4k)
frame_vm_group_bin_12643 = frame (4k)
frame_vm_group_bin_12644 = frame (4k)
frame_vm_group_bin_12645 = frame (4k)
frame_vm_group_bin_12646 = frame (4k)
frame_vm_group_bin_12647 = frame (4k)
frame_vm_group_bin_12648 = frame (4k)
frame_vm_group_bin_12649 = frame (4k)
frame_vm_group_bin_1265 = frame (4k)
frame_vm_group_bin_12650 = frame (4k)
frame_vm_group_bin_12651 = frame (4k)
frame_vm_group_bin_12652 = frame (4k)
frame_vm_group_bin_12653 = frame (4k)
frame_vm_group_bin_12654 = frame (4k)
frame_vm_group_bin_12655 = frame (4k)
frame_vm_group_bin_12656 = frame (4k)
frame_vm_group_bin_12657 = frame (4k)
frame_vm_group_bin_12658 = frame (4k)
frame_vm_group_bin_12659 = frame (4k)
frame_vm_group_bin_1266 = frame (4k)
frame_vm_group_bin_12660 = frame (4k)
frame_vm_group_bin_12661 = frame (4k)
frame_vm_group_bin_12662 = frame (4k)
frame_vm_group_bin_12663 = frame (4k)
frame_vm_group_bin_12664 = frame (4k)
frame_vm_group_bin_12665 = frame (4k)
frame_vm_group_bin_12666 = frame (4k)
frame_vm_group_bin_12667 = frame (4k)
frame_vm_group_bin_12668 = frame (4k)
frame_vm_group_bin_12669 = frame (4k)
frame_vm_group_bin_1267 = frame (4k)
frame_vm_group_bin_12670 = frame (4k)
frame_vm_group_bin_12671 = frame (4k)
frame_vm_group_bin_12672 = frame (4k)
frame_vm_group_bin_12673 = frame (4k)
frame_vm_group_bin_12674 = frame (4k)
frame_vm_group_bin_12675 = frame (4k)
frame_vm_group_bin_12676 = frame (4k)
frame_vm_group_bin_12677 = frame (4k)
frame_vm_group_bin_12678 = frame (4k)
frame_vm_group_bin_12679 = frame (4k)
frame_vm_group_bin_1268 = frame (4k)
frame_vm_group_bin_12680 = frame (4k)
frame_vm_group_bin_12681 = frame (4k)
frame_vm_group_bin_12682 = frame (4k)
frame_vm_group_bin_12683 = frame (4k)
frame_vm_group_bin_12684 = frame (4k)
frame_vm_group_bin_12685 = frame (4k)
frame_vm_group_bin_12686 = frame (4k)
frame_vm_group_bin_12687 = frame (4k)
frame_vm_group_bin_12688 = frame (4k)
frame_vm_group_bin_12689 = frame (4k)
frame_vm_group_bin_1269 = frame (4k)
frame_vm_group_bin_12690 = frame (4k)
frame_vm_group_bin_12691 = frame (4k)
frame_vm_group_bin_12692 = frame (4k)
frame_vm_group_bin_12693 = frame (4k)
frame_vm_group_bin_12694 = frame (4k)
frame_vm_group_bin_12695 = frame (4k)
frame_vm_group_bin_12696 = frame (4k)
frame_vm_group_bin_12697 = frame (4k)
frame_vm_group_bin_12698 = frame (4k)
frame_vm_group_bin_12699 = frame (4k)
frame_vm_group_bin_1270 = frame (4k)
frame_vm_group_bin_12700 = frame (4k)
frame_vm_group_bin_12701 = frame (4k)
frame_vm_group_bin_12702 = frame (4k)
frame_vm_group_bin_12703 = frame (4k)
frame_vm_group_bin_12704 = frame (4k)
frame_vm_group_bin_12705 = frame (4k)
frame_vm_group_bin_12706 = frame (4k)
frame_vm_group_bin_12707 = frame (4k)
frame_vm_group_bin_12708 = frame (4k)
frame_vm_group_bin_12709 = frame (4k)
frame_vm_group_bin_1271 = frame (4k)
frame_vm_group_bin_12710 = frame (4k)
frame_vm_group_bin_12711 = frame (4k)
frame_vm_group_bin_12712 = frame (4k)
frame_vm_group_bin_12713 = frame (4k)
frame_vm_group_bin_12714 = frame (4k)
frame_vm_group_bin_12715 = frame (4k)
frame_vm_group_bin_12716 = frame (4k)
frame_vm_group_bin_12717 = frame (4k)
frame_vm_group_bin_12718 = frame (4k)
frame_vm_group_bin_12719 = frame (4k)
frame_vm_group_bin_1272 = frame (4k)
frame_vm_group_bin_12720 = frame (4k)
frame_vm_group_bin_12721 = frame (4k)
frame_vm_group_bin_12722 = frame (4k)
frame_vm_group_bin_12723 = frame (4k)
frame_vm_group_bin_12724 = frame (4k)
frame_vm_group_bin_12725 = frame (4k)
frame_vm_group_bin_12726 = frame (4k)
frame_vm_group_bin_12727 = frame (4k)
frame_vm_group_bin_12728 = frame (4k)
frame_vm_group_bin_12729 = frame (4k)
frame_vm_group_bin_1273 = frame (4k)
frame_vm_group_bin_12730 = frame (4k)
frame_vm_group_bin_12731 = frame (4k)
frame_vm_group_bin_12732 = frame (4k)
frame_vm_group_bin_12733 = frame (4k)
frame_vm_group_bin_12734 = frame (4k)
frame_vm_group_bin_12735 = frame (4k)
frame_vm_group_bin_12736 = frame (4k)
frame_vm_group_bin_12737 = frame (4k)
frame_vm_group_bin_12738 = frame (4k)
frame_vm_group_bin_12739 = frame (4k)
frame_vm_group_bin_1274 = frame (4k)
frame_vm_group_bin_12740 = frame (4k)
frame_vm_group_bin_12741 = frame (4k)
frame_vm_group_bin_12742 = frame (4k)
frame_vm_group_bin_12743 = frame (4k)
frame_vm_group_bin_12744 = frame (4k)
frame_vm_group_bin_12745 = frame (4k)
frame_vm_group_bin_12746 = frame (4k)
frame_vm_group_bin_12747 = frame (4k)
frame_vm_group_bin_12748 = frame (4k)
frame_vm_group_bin_12749 = frame (4k)
frame_vm_group_bin_1275 = frame (4k)
frame_vm_group_bin_12750 = frame (4k)
frame_vm_group_bin_12751 = frame (4k)
frame_vm_group_bin_12752 = frame (4k)
frame_vm_group_bin_12753 = frame (4k)
frame_vm_group_bin_12754 = frame (4k)
frame_vm_group_bin_12755 = frame (4k)
frame_vm_group_bin_12756 = frame (4k)
frame_vm_group_bin_12757 = frame (4k)
frame_vm_group_bin_12758 = frame (4k)
frame_vm_group_bin_12759 = frame (4k)
frame_vm_group_bin_1276 = frame (4k)
frame_vm_group_bin_12760 = frame (4k)
frame_vm_group_bin_12761 = frame (4k)
frame_vm_group_bin_12762 = frame (4k)
frame_vm_group_bin_12763 = frame (4k)
frame_vm_group_bin_12764 = frame (4k)
frame_vm_group_bin_12765 = frame (4k)
frame_vm_group_bin_12766 = frame (4k)
frame_vm_group_bin_12767 = frame (4k)
frame_vm_group_bin_12768 = frame (4k)
frame_vm_group_bin_12769 = frame (4k)
frame_vm_group_bin_1277 = frame (4k)
frame_vm_group_bin_12770 = frame (4k)
frame_vm_group_bin_12771 = frame (4k)
frame_vm_group_bin_12772 = frame (4k)
frame_vm_group_bin_12773 = frame (4k)
frame_vm_group_bin_12774 = frame (4k)
frame_vm_group_bin_12775 = frame (4k)
frame_vm_group_bin_12776 = frame (4k)
frame_vm_group_bin_12777 = frame (4k)
frame_vm_group_bin_12778 = frame (4k)
frame_vm_group_bin_12779 = frame (4k)
frame_vm_group_bin_1278 = frame (4k)
frame_vm_group_bin_12780 = frame (4k)
frame_vm_group_bin_12781 = frame (4k)
frame_vm_group_bin_12782 = frame (4k)
frame_vm_group_bin_12783 = frame (4k)
frame_vm_group_bin_12784 = frame (4k)
frame_vm_group_bin_12785 = frame (4k)
frame_vm_group_bin_12786 = frame (4k)
frame_vm_group_bin_12787 = frame (4k)
frame_vm_group_bin_12788 = frame (4k)
frame_vm_group_bin_12789 = frame (4k)
frame_vm_group_bin_1279 = frame (4k)
frame_vm_group_bin_12790 = frame (4k)
frame_vm_group_bin_12791 = frame (4k)
frame_vm_group_bin_12792 = frame (4k)
frame_vm_group_bin_12793 = frame (4k)
frame_vm_group_bin_12794 = frame (4k)
frame_vm_group_bin_12795 = frame (4k)
frame_vm_group_bin_12796 = frame (4k)
frame_vm_group_bin_12797 = frame (4k)
frame_vm_group_bin_12798 = frame (4k)
frame_vm_group_bin_12799 = frame (4k)
frame_vm_group_bin_1280 = frame (4k)
frame_vm_group_bin_12800 = frame (4k)
frame_vm_group_bin_12801 = frame (4k)
frame_vm_group_bin_12802 = frame (4k)
frame_vm_group_bin_12803 = frame (4k)
frame_vm_group_bin_12804 = frame (4k)
frame_vm_group_bin_12805 = frame (4k)
frame_vm_group_bin_12806 = frame (4k)
frame_vm_group_bin_12807 = frame (4k)
frame_vm_group_bin_12808 = frame (4k)
frame_vm_group_bin_12809 = frame (4k)
frame_vm_group_bin_1281 = frame (4k)
frame_vm_group_bin_12810 = frame (4k)
frame_vm_group_bin_12811 = frame (4k)
frame_vm_group_bin_12812 = frame (4k)
frame_vm_group_bin_12813 = frame (4k)
frame_vm_group_bin_12814 = frame (4k)
frame_vm_group_bin_12815 = frame (4k)
frame_vm_group_bin_12816 = frame (4k)
frame_vm_group_bin_12817 = frame (4k)
frame_vm_group_bin_12818 = frame (4k)
frame_vm_group_bin_12819 = frame (4k)
frame_vm_group_bin_1282 = frame (4k)
frame_vm_group_bin_12820 = frame (4k)
frame_vm_group_bin_12821 = frame (4k)
frame_vm_group_bin_12822 = frame (4k)
frame_vm_group_bin_12823 = frame (4k)
frame_vm_group_bin_12824 = frame (4k)
frame_vm_group_bin_12825 = frame (4k)
frame_vm_group_bin_12826 = frame (4k)
frame_vm_group_bin_12827 = frame (4k)
frame_vm_group_bin_12828 = frame (4k)
frame_vm_group_bin_12829 = frame (4k)
frame_vm_group_bin_1283 = frame (4k)
frame_vm_group_bin_12830 = frame (4k)
frame_vm_group_bin_12831 = frame (4k)
frame_vm_group_bin_12832 = frame (4k)
frame_vm_group_bin_12833 = frame (4k)
frame_vm_group_bin_12834 = frame (4k)
frame_vm_group_bin_12835 = frame (4k)
frame_vm_group_bin_12836 = frame (4k)
frame_vm_group_bin_12837 = frame (4k)
frame_vm_group_bin_12838 = frame (4k)
frame_vm_group_bin_12839 = frame (4k)
frame_vm_group_bin_1284 = frame (4k)
frame_vm_group_bin_12840 = frame (4k)
frame_vm_group_bin_12841 = frame (4k)
frame_vm_group_bin_12842 = frame (4k)
frame_vm_group_bin_12843 = frame (4k)
frame_vm_group_bin_12844 = frame (4k)
frame_vm_group_bin_12845 = frame (4k)
frame_vm_group_bin_12846 = frame (4k)
frame_vm_group_bin_12847 = frame (4k)
frame_vm_group_bin_12848 = frame (4k)
frame_vm_group_bin_12849 = frame (4k)
frame_vm_group_bin_1285 = frame (4k)
frame_vm_group_bin_12850 = frame (4k)
frame_vm_group_bin_12851 = frame (4k)
frame_vm_group_bin_12852 = frame (4k)
frame_vm_group_bin_12853 = frame (4k)
frame_vm_group_bin_12854 = frame (4k)
frame_vm_group_bin_12855 = frame (4k)
frame_vm_group_bin_12856 = frame (4k)
frame_vm_group_bin_12857 = frame (4k)
frame_vm_group_bin_12858 = frame (4k)
frame_vm_group_bin_12859 = frame (4k)
frame_vm_group_bin_1286 = frame (4k)
frame_vm_group_bin_12860 = frame (4k)
frame_vm_group_bin_12861 = frame (4k)
frame_vm_group_bin_12862 = frame (4k)
frame_vm_group_bin_12863 = frame (4k)
frame_vm_group_bin_12864 = frame (4k)
frame_vm_group_bin_12865 = frame (4k)
frame_vm_group_bin_12866 = frame (4k)
frame_vm_group_bin_12867 = frame (4k)
frame_vm_group_bin_12868 = frame (4k)
frame_vm_group_bin_12869 = frame (4k)
frame_vm_group_bin_1287 = frame (4k)
frame_vm_group_bin_12870 = frame (4k)
frame_vm_group_bin_12871 = frame (4k)
frame_vm_group_bin_12872 = frame (4k)
frame_vm_group_bin_12873 = frame (4k)
frame_vm_group_bin_12874 = frame (4k)
frame_vm_group_bin_12875 = frame (4k)
frame_vm_group_bin_12876 = frame (4k)
frame_vm_group_bin_12877 = frame (4k)
frame_vm_group_bin_12878 = frame (4k)
frame_vm_group_bin_12879 = frame (4k)
frame_vm_group_bin_1288 = frame (4k)
frame_vm_group_bin_12880 = frame (4k)
frame_vm_group_bin_12881 = frame (4k)
frame_vm_group_bin_12882 = frame (4k)
frame_vm_group_bin_12883 = frame (4k)
frame_vm_group_bin_12884 = frame (4k)
frame_vm_group_bin_12885 = frame (4k)
frame_vm_group_bin_12886 = frame (4k)
frame_vm_group_bin_12887 = frame (4k)
frame_vm_group_bin_12888 = frame (4k)
frame_vm_group_bin_12889 = frame (4k)
frame_vm_group_bin_1289 = frame (4k)
frame_vm_group_bin_12890 = frame (4k)
frame_vm_group_bin_12891 = frame (4k)
frame_vm_group_bin_12892 = frame (4k)
frame_vm_group_bin_12893 = frame (4k)
frame_vm_group_bin_12894 = frame (4k)
frame_vm_group_bin_12895 = frame (4k)
frame_vm_group_bin_12896 = frame (4k)
frame_vm_group_bin_12897 = frame (4k)
frame_vm_group_bin_12898 = frame (4k)
frame_vm_group_bin_12899 = frame (4k)
frame_vm_group_bin_1290 = frame (4k)
frame_vm_group_bin_12900 = frame (4k)
frame_vm_group_bin_12901 = frame (4k)
frame_vm_group_bin_12902 = frame (4k)
frame_vm_group_bin_12903 = frame (4k)
frame_vm_group_bin_12904 = frame (4k)
frame_vm_group_bin_12905 = frame (4k)
frame_vm_group_bin_12906 = frame (4k)
frame_vm_group_bin_12907 = frame (4k)
frame_vm_group_bin_12908 = frame (4k)
frame_vm_group_bin_12909 = frame (4k)
frame_vm_group_bin_1291 = frame (4k)
frame_vm_group_bin_12910 = frame (4k)
frame_vm_group_bin_12911 = frame (4k)
frame_vm_group_bin_12912 = frame (4k)
frame_vm_group_bin_12913 = frame (4k)
frame_vm_group_bin_12914 = frame (4k)
frame_vm_group_bin_12915 = frame (4k)
frame_vm_group_bin_12916 = frame (4k)
frame_vm_group_bin_12917 = frame (4k)
frame_vm_group_bin_12918 = frame (4k)
frame_vm_group_bin_12919 = frame (4k)
frame_vm_group_bin_1292 = frame (4k)
frame_vm_group_bin_12920 = frame (4k)
frame_vm_group_bin_12921 = frame (4k)
frame_vm_group_bin_12922 = frame (4k)
frame_vm_group_bin_12923 = frame (4k)
frame_vm_group_bin_12924 = frame (4k)
frame_vm_group_bin_12925 = frame (4k)
frame_vm_group_bin_12926 = frame (4k)
frame_vm_group_bin_12927 = frame (4k)
frame_vm_group_bin_12928 = frame (4k)
frame_vm_group_bin_12929 = frame (4k)
frame_vm_group_bin_1293 = frame (4k)
frame_vm_group_bin_12930 = frame (4k)
frame_vm_group_bin_12931 = frame (4k)
frame_vm_group_bin_12932 = frame (4k)
frame_vm_group_bin_12933 = frame (4k)
frame_vm_group_bin_12934 = frame (4k)
frame_vm_group_bin_12935 = frame (4k)
frame_vm_group_bin_12936 = frame (4k)
frame_vm_group_bin_12937 = frame (4k)
frame_vm_group_bin_12938 = frame (4k)
frame_vm_group_bin_12939 = frame (4k)
frame_vm_group_bin_1294 = frame (4k)
frame_vm_group_bin_12940 = frame (4k)
frame_vm_group_bin_12941 = frame (4k)
frame_vm_group_bin_12942 = frame (4k)
frame_vm_group_bin_12943 = frame (4k)
frame_vm_group_bin_12944 = frame (4k)
frame_vm_group_bin_12945 = frame (4k)
frame_vm_group_bin_12946 = frame (4k)
frame_vm_group_bin_12947 = frame (4k)
frame_vm_group_bin_12948 = frame (4k)
frame_vm_group_bin_12949 = frame (4k)
frame_vm_group_bin_1295 = frame (4k)
frame_vm_group_bin_12950 = frame (4k)
frame_vm_group_bin_12951 = frame (4k)
frame_vm_group_bin_12952 = frame (4k)
frame_vm_group_bin_12953 = frame (4k)
frame_vm_group_bin_12954 = frame (4k)
frame_vm_group_bin_12955 = frame (4k)
frame_vm_group_bin_12956 = frame (4k)
frame_vm_group_bin_12957 = frame (4k)
frame_vm_group_bin_12958 = frame (4k)
frame_vm_group_bin_12959 = frame (4k)
frame_vm_group_bin_1296 = frame (4k)
frame_vm_group_bin_12960 = frame (4k)
frame_vm_group_bin_12961 = frame (4k)
frame_vm_group_bin_12962 = frame (4k)
frame_vm_group_bin_12963 = frame (4k)
frame_vm_group_bin_12964 = frame (4k)
frame_vm_group_bin_12965 = frame (4k)
frame_vm_group_bin_12966 = frame (4k)
frame_vm_group_bin_12967 = frame (4k)
frame_vm_group_bin_12968 = frame (4k)
frame_vm_group_bin_12969 = frame (4k)
frame_vm_group_bin_1297 = frame (4k)
frame_vm_group_bin_12970 = frame (4k)
frame_vm_group_bin_12971 = frame (4k)
frame_vm_group_bin_12972 = frame (4k)
frame_vm_group_bin_12973 = frame (4k)
frame_vm_group_bin_12974 = frame (4k)
frame_vm_group_bin_12975 = frame (4k)
frame_vm_group_bin_12976 = frame (4k)
frame_vm_group_bin_12977 = frame (4k)
frame_vm_group_bin_12978 = frame (4k)
frame_vm_group_bin_12979 = frame (4k)
frame_vm_group_bin_1298 = frame (4k)
frame_vm_group_bin_12980 = frame (4k)
frame_vm_group_bin_12981 = frame (4k)
frame_vm_group_bin_12982 = frame (4k)
frame_vm_group_bin_12983 = frame (4k)
frame_vm_group_bin_12984 = frame (4k)
frame_vm_group_bin_12985 = frame (4k)
frame_vm_group_bin_12986 = frame (4k)
frame_vm_group_bin_12987 = frame (4k)
frame_vm_group_bin_12988 = frame (4k)
frame_vm_group_bin_12989 = frame (4k)
frame_vm_group_bin_1299 = frame (4k)
frame_vm_group_bin_12990 = frame (4k)
frame_vm_group_bin_12991 = frame (4k)
frame_vm_group_bin_12992 = frame (4k)
frame_vm_group_bin_12993 = frame (4k)
frame_vm_group_bin_12994 = frame (4k)
frame_vm_group_bin_12995 = frame (4k)
frame_vm_group_bin_12996 = frame (4k)
frame_vm_group_bin_12997 = frame (4k)
frame_vm_group_bin_12998 = frame (4k)
frame_vm_group_bin_12999 = frame (4k)
frame_vm_group_bin_1300 = frame (4k)
frame_vm_group_bin_13000 = frame (4k)
frame_vm_group_bin_13001 = frame (4k)
frame_vm_group_bin_13002 = frame (4k)
frame_vm_group_bin_13003 = frame (4k)
frame_vm_group_bin_13004 = frame (4k)
frame_vm_group_bin_13005 = frame (4k)
frame_vm_group_bin_13006 = frame (4k)
frame_vm_group_bin_13007 = frame (4k)
frame_vm_group_bin_13008 = frame (4k)
frame_vm_group_bin_13009 = frame (4k)
frame_vm_group_bin_1301 = frame (4k)
frame_vm_group_bin_13010 = frame (4k)
frame_vm_group_bin_13011 = frame (4k)
frame_vm_group_bin_13012 = frame (4k)
frame_vm_group_bin_13013 = frame (4k)
frame_vm_group_bin_13014 = frame (4k)
frame_vm_group_bin_13015 = frame (4k)
frame_vm_group_bin_13016 = frame (4k)
frame_vm_group_bin_13017 = frame (4k)
frame_vm_group_bin_13018 = frame (4k)
frame_vm_group_bin_13019 = frame (4k)
frame_vm_group_bin_1302 = frame (4k)
frame_vm_group_bin_13020 = frame (4k)
frame_vm_group_bin_13021 = frame (4k)
frame_vm_group_bin_13022 = frame (4k)
frame_vm_group_bin_13023 = frame (4k)
frame_vm_group_bin_13024 = frame (4k)
frame_vm_group_bin_13025 = frame (4k)
frame_vm_group_bin_13026 = frame (4k)
frame_vm_group_bin_13027 = frame (4k)
frame_vm_group_bin_13028 = frame (4k)
frame_vm_group_bin_13029 = frame (4k)
frame_vm_group_bin_1303 = frame (4k)
frame_vm_group_bin_13030 = frame (4k)
frame_vm_group_bin_13031 = frame (4k)
frame_vm_group_bin_13032 = frame (4k)
frame_vm_group_bin_13033 = frame (4k)
frame_vm_group_bin_13034 = frame (4k)
frame_vm_group_bin_13035 = frame (4k)
frame_vm_group_bin_13036 = frame (4k)
frame_vm_group_bin_13037 = frame (4k)
frame_vm_group_bin_13038 = frame (4k)
frame_vm_group_bin_13039 = frame (4k)
frame_vm_group_bin_1304 = frame (4k)
frame_vm_group_bin_13040 = frame (4k)
frame_vm_group_bin_13041 = frame (4k)
frame_vm_group_bin_13042 = frame (4k)
frame_vm_group_bin_13043 = frame (4k)
frame_vm_group_bin_13044 = frame (4k)
frame_vm_group_bin_13045 = frame (4k)
frame_vm_group_bin_13046 = frame (4k)
frame_vm_group_bin_13047 = frame (4k)
frame_vm_group_bin_13048 = frame (4k)
frame_vm_group_bin_13049 = frame (4k)
frame_vm_group_bin_1305 = frame (4k)
frame_vm_group_bin_13050 = frame (4k)
frame_vm_group_bin_13051 = frame (4k)
frame_vm_group_bin_13052 = frame (4k)
frame_vm_group_bin_13053 = frame (4k)
frame_vm_group_bin_13054 = frame (4k)
frame_vm_group_bin_13055 = frame (4k)
frame_vm_group_bin_13056 = frame (4k)
frame_vm_group_bin_13057 = frame (4k)
frame_vm_group_bin_13058 = frame (4k)
frame_vm_group_bin_13059 = frame (4k)
frame_vm_group_bin_1306 = frame (4k)
frame_vm_group_bin_13060 = frame (4k)
frame_vm_group_bin_13061 = frame (4k)
frame_vm_group_bin_13062 = frame (4k)
frame_vm_group_bin_13063 = frame (4k)
frame_vm_group_bin_13064 = frame (4k)
frame_vm_group_bin_13065 = frame (4k)
frame_vm_group_bin_13066 = frame (4k)
frame_vm_group_bin_13067 = frame (4k)
frame_vm_group_bin_13068 = frame (4k)
frame_vm_group_bin_13069 = frame (4k)
frame_vm_group_bin_1307 = frame (4k)
frame_vm_group_bin_13070 = frame (4k)
frame_vm_group_bin_13071 = frame (4k)
frame_vm_group_bin_13072 = frame (4k)
frame_vm_group_bin_13073 = frame (4k)
frame_vm_group_bin_13074 = frame (4k)
frame_vm_group_bin_13075 = frame (4k)
frame_vm_group_bin_13076 = frame (4k)
frame_vm_group_bin_13077 = frame (4k)
frame_vm_group_bin_13078 = frame (4k)
frame_vm_group_bin_13079 = frame (4k)
frame_vm_group_bin_1308 = frame (4k)
frame_vm_group_bin_13080 = frame (4k)
frame_vm_group_bin_13081 = frame (4k)
frame_vm_group_bin_13082 = frame (4k)
frame_vm_group_bin_13083 = frame (4k)
frame_vm_group_bin_13084 = frame (4k)
frame_vm_group_bin_13085 = frame (4k)
frame_vm_group_bin_13086 = frame (4k)
frame_vm_group_bin_13087 = frame (4k)
frame_vm_group_bin_13088 = frame (4k)
frame_vm_group_bin_13089 = frame (4k)
frame_vm_group_bin_1309 = frame (4k)
frame_vm_group_bin_13090 = frame (4k)
frame_vm_group_bin_13091 = frame (4k)
frame_vm_group_bin_13092 = frame (4k)
frame_vm_group_bin_13093 = frame (4k)
frame_vm_group_bin_13094 = frame (4k)
frame_vm_group_bin_13095 = frame (4k)
frame_vm_group_bin_13096 = frame (4k)
frame_vm_group_bin_13097 = frame (4k)
frame_vm_group_bin_13098 = frame (4k)
frame_vm_group_bin_13099 = frame (4k)
frame_vm_group_bin_1310 = frame (4k)
frame_vm_group_bin_13100 = frame (4k)
frame_vm_group_bin_13101 = frame (4k)
frame_vm_group_bin_13102 = frame (4k)
frame_vm_group_bin_13103 = frame (4k)
frame_vm_group_bin_13104 = frame (4k)
frame_vm_group_bin_13105 = frame (4k)
frame_vm_group_bin_13106 = frame (4k)
frame_vm_group_bin_13107 = frame (4k)
frame_vm_group_bin_13108 = frame (4k)
frame_vm_group_bin_13109 = frame (4k)
frame_vm_group_bin_1311 = frame (4k)
frame_vm_group_bin_13110 = frame (4k)
frame_vm_group_bin_13111 = frame (4k)
frame_vm_group_bin_13112 = frame (4k)
frame_vm_group_bin_13113 = frame (4k)
frame_vm_group_bin_13114 = frame (4k)
frame_vm_group_bin_13115 = frame (4k)
frame_vm_group_bin_13116 = frame (4k)
frame_vm_group_bin_13117 = frame (4k)
frame_vm_group_bin_13118 = frame (4k)
frame_vm_group_bin_13119 = frame (4k)
frame_vm_group_bin_1312 = frame (4k)
frame_vm_group_bin_13120 = frame (4k)
frame_vm_group_bin_13121 = frame (4k)
frame_vm_group_bin_13122 = frame (4k)
frame_vm_group_bin_13123 = frame (4k)
frame_vm_group_bin_13124 = frame (4k)
frame_vm_group_bin_13125 = frame (4k)
frame_vm_group_bin_13126 = frame (4k)
frame_vm_group_bin_13127 = frame (4k)
frame_vm_group_bin_13128 = frame (4k)
frame_vm_group_bin_13129 = frame (4k)
frame_vm_group_bin_1313 = frame (4k)
frame_vm_group_bin_13130 = frame (4k)
frame_vm_group_bin_13131 = frame (4k)
frame_vm_group_bin_13132 = frame (4k)
frame_vm_group_bin_13133 = frame (4k)
frame_vm_group_bin_13134 = frame (4k)
frame_vm_group_bin_13135 = frame (4k)
frame_vm_group_bin_13136 = frame (4k)
frame_vm_group_bin_13137 = frame (4k)
frame_vm_group_bin_13138 = frame (4k)
frame_vm_group_bin_13139 = frame (4k)
frame_vm_group_bin_1314 = frame (4k)
frame_vm_group_bin_13140 = frame (4k)
frame_vm_group_bin_13141 = frame (4k)
frame_vm_group_bin_13142 = frame (4k)
frame_vm_group_bin_13143 = frame (4k)
frame_vm_group_bin_13144 = frame (4k)
frame_vm_group_bin_13145 = frame (4k)
frame_vm_group_bin_13146 = frame (4k)
frame_vm_group_bin_13147 = frame (4k)
frame_vm_group_bin_13148 = frame (4k)
frame_vm_group_bin_13149 = frame (4k)
frame_vm_group_bin_1315 = frame (4k)
frame_vm_group_bin_13150 = frame (4k)
frame_vm_group_bin_13151 = frame (4k)
frame_vm_group_bin_13152 = frame (4k)
frame_vm_group_bin_13153 = frame (4k)
frame_vm_group_bin_13154 = frame (4k)
frame_vm_group_bin_13155 = frame (4k)
frame_vm_group_bin_13156 = frame (4k)
frame_vm_group_bin_13157 = frame (4k)
frame_vm_group_bin_13158 = frame (4k)
frame_vm_group_bin_13159 = frame (4k)
frame_vm_group_bin_1316 = frame (4k)
frame_vm_group_bin_13160 = frame (4k)
frame_vm_group_bin_13161 = frame (4k)
frame_vm_group_bin_13162 = frame (4k)
frame_vm_group_bin_13163 = frame (4k)
frame_vm_group_bin_13164 = frame (4k)
frame_vm_group_bin_13165 = frame (4k)
frame_vm_group_bin_13166 = frame (4k)
frame_vm_group_bin_13167 = frame (4k)
frame_vm_group_bin_13168 = frame (4k)
frame_vm_group_bin_13169 = frame (4k)
frame_vm_group_bin_1317 = frame (4k)
frame_vm_group_bin_13170 = frame (4k)
frame_vm_group_bin_13171 = frame (4k)
frame_vm_group_bin_13172 = frame (4k)
frame_vm_group_bin_13173 = frame (4k)
frame_vm_group_bin_13174 = frame (4k)
frame_vm_group_bin_13175 = frame (4k)
frame_vm_group_bin_13176 = frame (4k)
frame_vm_group_bin_13177 = frame (4k)
frame_vm_group_bin_13178 = frame (4k)
frame_vm_group_bin_13179 = frame (4k)
frame_vm_group_bin_1318 = frame (4k)
frame_vm_group_bin_13180 = frame (4k)
frame_vm_group_bin_13181 = frame (4k)
frame_vm_group_bin_13182 = frame (4k)
frame_vm_group_bin_13183 = frame (4k)
frame_vm_group_bin_13184 = frame (4k)
frame_vm_group_bin_13185 = frame (4k)
frame_vm_group_bin_13186 = frame (4k)
frame_vm_group_bin_13187 = frame (4k)
frame_vm_group_bin_13188 = frame (4k)
frame_vm_group_bin_13189 = frame (4k)
frame_vm_group_bin_1319 = frame (4k)
frame_vm_group_bin_13190 = frame (4k)
frame_vm_group_bin_13191 = frame (4k)
frame_vm_group_bin_13192 = frame (4k)
frame_vm_group_bin_13193 = frame (4k)
frame_vm_group_bin_13194 = frame (4k)
frame_vm_group_bin_13195 = frame (4k)
frame_vm_group_bin_13196 = frame (4k)
frame_vm_group_bin_13197 = frame (4k)
frame_vm_group_bin_13198 = frame (4k)
frame_vm_group_bin_13199 = frame (4k)
frame_vm_group_bin_1320 = frame (4k)
frame_vm_group_bin_13200 = frame (4k)
frame_vm_group_bin_13201 = frame (4k)
frame_vm_group_bin_13202 = frame (4k)
frame_vm_group_bin_13203 = frame (4k)
frame_vm_group_bin_13204 = frame (4k)
frame_vm_group_bin_13205 = frame (4k)
frame_vm_group_bin_13206 = frame (4k)
frame_vm_group_bin_13207 = frame (4k)
frame_vm_group_bin_13208 = frame (4k)
frame_vm_group_bin_13209 = frame (4k)
frame_vm_group_bin_1321 = frame (4k)
frame_vm_group_bin_13210 = frame (4k)
frame_vm_group_bin_13211 = frame (4k)
frame_vm_group_bin_13212 = frame (4k)
frame_vm_group_bin_13213 = frame (4k)
frame_vm_group_bin_13214 = frame (4k)
frame_vm_group_bin_13215 = frame (4k)
frame_vm_group_bin_13216 = frame (4k)
frame_vm_group_bin_13217 = frame (4k)
frame_vm_group_bin_13218 = frame (4k)
frame_vm_group_bin_13219 = frame (4k)
frame_vm_group_bin_1322 = frame (4k)
frame_vm_group_bin_13220 = frame (4k)
frame_vm_group_bin_13221 = frame (4k)
frame_vm_group_bin_13222 = frame (4k)
frame_vm_group_bin_13223 = frame (4k)
frame_vm_group_bin_13224 = frame (4k)
frame_vm_group_bin_13225 = frame (4k)
frame_vm_group_bin_13226 = frame (4k)
frame_vm_group_bin_13227 = frame (4k)
frame_vm_group_bin_13228 = frame (4k)
frame_vm_group_bin_13229 = frame (4k)
frame_vm_group_bin_1323 = frame (4k)
frame_vm_group_bin_13230 = frame (4k)
frame_vm_group_bin_13231 = frame (4k)
frame_vm_group_bin_13232 = frame (4k)
frame_vm_group_bin_13233 = frame (4k)
frame_vm_group_bin_13234 = frame (4k)
frame_vm_group_bin_13235 = frame (4k)
frame_vm_group_bin_13236 = frame (4k)
frame_vm_group_bin_13237 = frame (4k)
frame_vm_group_bin_13238 = frame (4k)
frame_vm_group_bin_13239 = frame (4k)
frame_vm_group_bin_1324 = frame (4k)
frame_vm_group_bin_13240 = frame (4k)
frame_vm_group_bin_13241 = frame (4k)
frame_vm_group_bin_13242 = frame (4k)
frame_vm_group_bin_13243 = frame (4k)
frame_vm_group_bin_13244 = frame (4k)
frame_vm_group_bin_13245 = frame (4k)
frame_vm_group_bin_13246 = frame (4k)
frame_vm_group_bin_13247 = frame (4k)
frame_vm_group_bin_13248 = frame (4k)
frame_vm_group_bin_13249 = frame (4k)
frame_vm_group_bin_1325 = frame (4k)
frame_vm_group_bin_13250 = frame (4k)
frame_vm_group_bin_13251 = frame (4k)
frame_vm_group_bin_13252 = frame (4k)
frame_vm_group_bin_13253 = frame (4k)
frame_vm_group_bin_13254 = frame (4k)
frame_vm_group_bin_13255 = frame (4k)
frame_vm_group_bin_13256 = frame (4k)
frame_vm_group_bin_13257 = frame (4k)
frame_vm_group_bin_13258 = frame (4k)
frame_vm_group_bin_13259 = frame (4k)
frame_vm_group_bin_1326 = frame (4k)
frame_vm_group_bin_13260 = frame (4k)
frame_vm_group_bin_13261 = frame (4k)
frame_vm_group_bin_13262 = frame (4k)
frame_vm_group_bin_13263 = frame (4k)
frame_vm_group_bin_13264 = frame (4k)
frame_vm_group_bin_13265 = frame (4k)
frame_vm_group_bin_13266 = frame (4k)
frame_vm_group_bin_13267 = frame (4k)
frame_vm_group_bin_13268 = frame (4k)
frame_vm_group_bin_13269 = frame (4k)
frame_vm_group_bin_1327 = frame (4k)
frame_vm_group_bin_13270 = frame (4k)
frame_vm_group_bin_13271 = frame (4k)
frame_vm_group_bin_13272 = frame (4k)
frame_vm_group_bin_13273 = frame (4k)
frame_vm_group_bin_13274 = frame (4k)
frame_vm_group_bin_13275 = frame (4k)
frame_vm_group_bin_13276 = frame (4k)
frame_vm_group_bin_13277 = frame (4k)
frame_vm_group_bin_13278 = frame (4k)
frame_vm_group_bin_13279 = frame (4k)
frame_vm_group_bin_1328 = frame (4k)
frame_vm_group_bin_13280 = frame (4k)
frame_vm_group_bin_13281 = frame (4k)
frame_vm_group_bin_13282 = frame (4k)
frame_vm_group_bin_13283 = frame (4k)
frame_vm_group_bin_13284 = frame (4k)
frame_vm_group_bin_13285 = frame (4k)
frame_vm_group_bin_13286 = frame (4k)
frame_vm_group_bin_13287 = frame (4k)
frame_vm_group_bin_13288 = frame (4k)
frame_vm_group_bin_13289 = frame (4k)
frame_vm_group_bin_1329 = frame (4k)
frame_vm_group_bin_13290 = frame (4k)
frame_vm_group_bin_13291 = frame (4k)
frame_vm_group_bin_13292 = frame (4k)
frame_vm_group_bin_13293 = frame (4k)
frame_vm_group_bin_13294 = frame (4k)
frame_vm_group_bin_13295 = frame (4k)
frame_vm_group_bin_13296 = frame (4k)
frame_vm_group_bin_13297 = frame (4k)
frame_vm_group_bin_13298 = frame (4k)
frame_vm_group_bin_13299 = frame (4k)
frame_vm_group_bin_1330 = frame (4k)
frame_vm_group_bin_13300 = frame (4k)
frame_vm_group_bin_13301 = frame (4k)
frame_vm_group_bin_13302 = frame (4k)
frame_vm_group_bin_13303 = frame (4k)
frame_vm_group_bin_13304 = frame (4k)
frame_vm_group_bin_13305 = frame (4k)
frame_vm_group_bin_13306 = frame (4k)
frame_vm_group_bin_13307 = frame (4k)
frame_vm_group_bin_13308 = frame (4k)
frame_vm_group_bin_13309 = frame (4k)
frame_vm_group_bin_1331 = frame (4k)
frame_vm_group_bin_13310 = frame (4k)
frame_vm_group_bin_13311 = frame (4k)
frame_vm_group_bin_13312 = frame (4k)
frame_vm_group_bin_13313 = frame (4k)
frame_vm_group_bin_13314 = frame (4k)
frame_vm_group_bin_13315 = frame (4k)
frame_vm_group_bin_13316 = frame (4k)
frame_vm_group_bin_13317 = frame (4k)
frame_vm_group_bin_13318 = frame (4k)
frame_vm_group_bin_13319 = frame (4k)
frame_vm_group_bin_1332 = frame (4k)
frame_vm_group_bin_13320 = frame (4k)
frame_vm_group_bin_13321 = frame (4k)
frame_vm_group_bin_13322 = frame (4k)
frame_vm_group_bin_13323 = frame (4k)
frame_vm_group_bin_13324 = frame (4k)
frame_vm_group_bin_13325 = frame (4k)
frame_vm_group_bin_13326 = frame (4k)
frame_vm_group_bin_13327 = frame (4k)
frame_vm_group_bin_13328 = frame (4k)
frame_vm_group_bin_13329 = frame (4k)
frame_vm_group_bin_1333 = frame (4k)
frame_vm_group_bin_13330 = frame (4k)
frame_vm_group_bin_13331 = frame (4k)
frame_vm_group_bin_13332 = frame (4k)
frame_vm_group_bin_13333 = frame (4k)
frame_vm_group_bin_13334 = frame (4k)
frame_vm_group_bin_13335 = frame (4k)
frame_vm_group_bin_13336 = frame (4k)
frame_vm_group_bin_13337 = frame (4k)
frame_vm_group_bin_13338 = frame (4k)
frame_vm_group_bin_13339 = frame (4k)
frame_vm_group_bin_1334 = frame (4k)
frame_vm_group_bin_13340 = frame (4k)
frame_vm_group_bin_13341 = frame (4k)
frame_vm_group_bin_13342 = frame (4k)
frame_vm_group_bin_13343 = frame (4k)
frame_vm_group_bin_13344 = frame (4k)
frame_vm_group_bin_13345 = frame (4k)
frame_vm_group_bin_13346 = frame (4k)
frame_vm_group_bin_13347 = frame (4k)
frame_vm_group_bin_13348 = frame (4k)
frame_vm_group_bin_13349 = frame (4k)
frame_vm_group_bin_1335 = frame (4k)
frame_vm_group_bin_13350 = frame (4k)
frame_vm_group_bin_13351 = frame (4k)
frame_vm_group_bin_13352 = frame (4k)
frame_vm_group_bin_13353 = frame (4k)
frame_vm_group_bin_13354 = frame (4k)
frame_vm_group_bin_13355 = frame (4k)
frame_vm_group_bin_13356 = frame (4k)
frame_vm_group_bin_13357 = frame (4k)
frame_vm_group_bin_13358 = frame (4k)
frame_vm_group_bin_13359 = frame (4k)
frame_vm_group_bin_1336 = frame (4k)
frame_vm_group_bin_13360 = frame (4k)
frame_vm_group_bin_13361 = frame (4k)
frame_vm_group_bin_13362 = frame (4k)
frame_vm_group_bin_13363 = frame (4k)
frame_vm_group_bin_13364 = frame (4k)
frame_vm_group_bin_13365 = frame (4k)
frame_vm_group_bin_13366 = frame (4k)
frame_vm_group_bin_13367 = frame (4k)
frame_vm_group_bin_13368 = frame (4k)
frame_vm_group_bin_13369 = frame (4k)
frame_vm_group_bin_1337 = frame (4k)
frame_vm_group_bin_13370 = frame (4k)
frame_vm_group_bin_13371 = frame (4k)
frame_vm_group_bin_13372 = frame (4k)
frame_vm_group_bin_13373 = frame (4k)
frame_vm_group_bin_13374 = frame (4k)
frame_vm_group_bin_13375 = frame (4k)
frame_vm_group_bin_13376 = frame (4k)
frame_vm_group_bin_13377 = frame (4k)
frame_vm_group_bin_13378 = frame (4k)
frame_vm_group_bin_13379 = frame (4k)
frame_vm_group_bin_1338 = frame (4k)
frame_vm_group_bin_13380 = frame (4k)
frame_vm_group_bin_13381 = frame (4k)
frame_vm_group_bin_13382 = frame (4k)
frame_vm_group_bin_13383 = frame (4k)
frame_vm_group_bin_13384 = frame (4k)
frame_vm_group_bin_13385 = frame (4k)
frame_vm_group_bin_13386 = frame (4k)
frame_vm_group_bin_13387 = frame (4k)
frame_vm_group_bin_13388 = frame (4k)
frame_vm_group_bin_13389 = frame (4k)
frame_vm_group_bin_1339 = frame (4k)
frame_vm_group_bin_13390 = frame (4k)
frame_vm_group_bin_13391 = frame (4k)
frame_vm_group_bin_13392 = frame (4k)
frame_vm_group_bin_13393 = frame (4k)
frame_vm_group_bin_13394 = frame (4k)
frame_vm_group_bin_13395 = frame (4k)
frame_vm_group_bin_13396 = frame (4k)
frame_vm_group_bin_13397 = frame (4k)
frame_vm_group_bin_13398 = frame (4k)
frame_vm_group_bin_13399 = frame (4k)
frame_vm_group_bin_1340 = frame (4k)
frame_vm_group_bin_13400 = frame (4k)
frame_vm_group_bin_13401 = frame (4k)
frame_vm_group_bin_13402 = frame (4k)
frame_vm_group_bin_13403 = frame (4k)
frame_vm_group_bin_13404 = frame (4k)
frame_vm_group_bin_13405 = frame (4k)
frame_vm_group_bin_13406 = frame (4k)
frame_vm_group_bin_13407 = frame (4k)
frame_vm_group_bin_13408 = frame (4k)
frame_vm_group_bin_13409 = frame (4k)
frame_vm_group_bin_1341 = frame (4k)
frame_vm_group_bin_13410 = frame (4k)
frame_vm_group_bin_13411 = frame (4k)
frame_vm_group_bin_13412 = frame (4k)
frame_vm_group_bin_13413 = frame (4k)
frame_vm_group_bin_13414 = frame (4k)
frame_vm_group_bin_13415 = frame (4k)
frame_vm_group_bin_13416 = frame (4k)
frame_vm_group_bin_13417 = frame (4k)
frame_vm_group_bin_13418 = frame (4k)
frame_vm_group_bin_13419 = frame (4k)
frame_vm_group_bin_1342 = frame (4k)
frame_vm_group_bin_13420 = frame (4k)
frame_vm_group_bin_13421 = frame (4k)
frame_vm_group_bin_13422 = frame (4k)
frame_vm_group_bin_13423 = frame (4k)
frame_vm_group_bin_13424 = frame (4k)
frame_vm_group_bin_13425 = frame (4k)
frame_vm_group_bin_13426 = frame (4k)
frame_vm_group_bin_13427 = frame (4k)
frame_vm_group_bin_13428 = frame (4k)
frame_vm_group_bin_13429 = frame (4k)
frame_vm_group_bin_1343 = frame (4k)
frame_vm_group_bin_13430 = frame (4k)
frame_vm_group_bin_13431 = frame (4k)
frame_vm_group_bin_13432 = frame (4k)
frame_vm_group_bin_13433 = frame (4k)
frame_vm_group_bin_13434 = frame (4k)
frame_vm_group_bin_13435 = frame (4k)
frame_vm_group_bin_13436 = frame (4k)
frame_vm_group_bin_13437 = frame (4k)
frame_vm_group_bin_13438 = frame (4k)
frame_vm_group_bin_13439 = frame (4k)
frame_vm_group_bin_1344 = frame (4k)
frame_vm_group_bin_13440 = frame (4k)
frame_vm_group_bin_13441 = frame (4k)
frame_vm_group_bin_13442 = frame (4k)
frame_vm_group_bin_13443 = frame (4k)
frame_vm_group_bin_13444 = frame (4k)
frame_vm_group_bin_13445 = frame (4k)
frame_vm_group_bin_13446 = frame (4k)
frame_vm_group_bin_13447 = frame (4k)
frame_vm_group_bin_13448 = frame (4k)
frame_vm_group_bin_13449 = frame (4k)
frame_vm_group_bin_1345 = frame (4k)
frame_vm_group_bin_13450 = frame (4k)
frame_vm_group_bin_13451 = frame (4k)
frame_vm_group_bin_13452 = frame (4k)
frame_vm_group_bin_13453 = frame (4k)
frame_vm_group_bin_13454 = frame (4k)
frame_vm_group_bin_13455 = frame (4k)
frame_vm_group_bin_13456 = frame (4k)
frame_vm_group_bin_13457 = frame (4k)
frame_vm_group_bin_13458 = frame (4k)
frame_vm_group_bin_13459 = frame (4k)
frame_vm_group_bin_1346 = frame (4k)
frame_vm_group_bin_13460 = frame (4k)
frame_vm_group_bin_13461 = frame (4k)
frame_vm_group_bin_13462 = frame (4k)
frame_vm_group_bin_13463 = frame (4k)
frame_vm_group_bin_13464 = frame (4k)
frame_vm_group_bin_13465 = frame (4k)
frame_vm_group_bin_13466 = frame (4k)
frame_vm_group_bin_13467 = frame (4k)
frame_vm_group_bin_13468 = frame (4k)
frame_vm_group_bin_13469 = frame (4k)
frame_vm_group_bin_1347 = frame (4k)
frame_vm_group_bin_13470 = frame (4k)
frame_vm_group_bin_13471 = frame (4k)
frame_vm_group_bin_13472 = frame (4k)
frame_vm_group_bin_13473 = frame (4k)
frame_vm_group_bin_13474 = frame (4k)
frame_vm_group_bin_13475 = frame (4k)
frame_vm_group_bin_13476 = frame (4k)
frame_vm_group_bin_13477 = frame (4k)
frame_vm_group_bin_13478 = frame (4k)
frame_vm_group_bin_13479 = frame (4k)
frame_vm_group_bin_1348 = frame (4k)
frame_vm_group_bin_13480 = frame (4k)
frame_vm_group_bin_13481 = frame (4k)
frame_vm_group_bin_13482 = frame (4k)
frame_vm_group_bin_13483 = frame (4k)
frame_vm_group_bin_13484 = frame (4k)
frame_vm_group_bin_13485 = frame (4k)
frame_vm_group_bin_13486 = frame (4k)
frame_vm_group_bin_13487 = frame (4k)
frame_vm_group_bin_13488 = frame (4k)
frame_vm_group_bin_13489 = frame (4k)
frame_vm_group_bin_1349 = frame (4k)
frame_vm_group_bin_13490 = frame (4k)
frame_vm_group_bin_13491 = frame (4k)
frame_vm_group_bin_13492 = frame (4k)
frame_vm_group_bin_13493 = frame (4k)
frame_vm_group_bin_13494 = frame (4k)
frame_vm_group_bin_13495 = frame (4k)
frame_vm_group_bin_13496 = frame (4k)
frame_vm_group_bin_13497 = frame (4k)
frame_vm_group_bin_13498 = frame (4k)
frame_vm_group_bin_13499 = frame (4k)
frame_vm_group_bin_1350 = frame (4k)
frame_vm_group_bin_13500 = frame (4k)
frame_vm_group_bin_13501 = frame (4k)
frame_vm_group_bin_13502 = frame (4k)
frame_vm_group_bin_13503 = frame (4k)
frame_vm_group_bin_13504 = frame (4k)
frame_vm_group_bin_13505 = frame (4k)
frame_vm_group_bin_13506 = frame (4k)
frame_vm_group_bin_13507 = frame (4k)
frame_vm_group_bin_13508 = frame (4k)
frame_vm_group_bin_13509 = frame (4k)
frame_vm_group_bin_1351 = frame (4k)
frame_vm_group_bin_13510 = frame (4k)
frame_vm_group_bin_13511 = frame (4k)
frame_vm_group_bin_13512 = frame (4k)
frame_vm_group_bin_13513 = frame (4k)
frame_vm_group_bin_13514 = frame (4k)
frame_vm_group_bin_13515 = frame (4k)
frame_vm_group_bin_13516 = frame (4k)
frame_vm_group_bin_13517 = frame (4k)
frame_vm_group_bin_13518 = frame (4k)
frame_vm_group_bin_13519 = frame (4k)
frame_vm_group_bin_1352 = frame (4k)
frame_vm_group_bin_13520 = frame (4k)
frame_vm_group_bin_13521 = frame (4k)
frame_vm_group_bin_13522 = frame (4k)
frame_vm_group_bin_13523 = frame (4k)
frame_vm_group_bin_13524 = frame (4k)
frame_vm_group_bin_13525 = frame (4k)
frame_vm_group_bin_13526 = frame (4k)
frame_vm_group_bin_13527 = frame (4k)
frame_vm_group_bin_13528 = frame (4k)
frame_vm_group_bin_13529 = frame (4k)
frame_vm_group_bin_1353 = frame (4k)
frame_vm_group_bin_13530 = frame (4k)
frame_vm_group_bin_13531 = frame (4k)
frame_vm_group_bin_13532 = frame (4k)
frame_vm_group_bin_13533 = frame (4k)
frame_vm_group_bin_13534 = frame (4k)
frame_vm_group_bin_13535 = frame (4k)
frame_vm_group_bin_13536 = frame (4k)
frame_vm_group_bin_13537 = frame (4k)
frame_vm_group_bin_13538 = frame (4k)
frame_vm_group_bin_13539 = frame (4k)
frame_vm_group_bin_1354 = frame (4k)
frame_vm_group_bin_13540 = frame (4k)
frame_vm_group_bin_13541 = frame (4k)
frame_vm_group_bin_13542 = frame (4k)
frame_vm_group_bin_13543 = frame (4k)
frame_vm_group_bin_13544 = frame (4k)
frame_vm_group_bin_13545 = frame (4k)
frame_vm_group_bin_13546 = frame (4k)
frame_vm_group_bin_13547 = frame (4k)
frame_vm_group_bin_13548 = frame (4k)
frame_vm_group_bin_13549 = frame (4k)
frame_vm_group_bin_1355 = frame (4k)
frame_vm_group_bin_13550 = frame (4k)
frame_vm_group_bin_13551 = frame (4k)
frame_vm_group_bin_13552 = frame (4k)
frame_vm_group_bin_13553 = frame (4k)
frame_vm_group_bin_13554 = frame (4k)
frame_vm_group_bin_13555 = frame (4k)
frame_vm_group_bin_13556 = frame (4k)
frame_vm_group_bin_13557 = frame (4k)
frame_vm_group_bin_13558 = frame (4k)
frame_vm_group_bin_13559 = frame (4k)
frame_vm_group_bin_1356 = frame (4k)
frame_vm_group_bin_13560 = frame (4k)
frame_vm_group_bin_13561 = frame (4k)
frame_vm_group_bin_13562 = frame (4k)
frame_vm_group_bin_13563 = frame (4k)
frame_vm_group_bin_13564 = frame (4k)
frame_vm_group_bin_13565 = frame (4k)
frame_vm_group_bin_13566 = frame (4k)
frame_vm_group_bin_13567 = frame (4k)
frame_vm_group_bin_13568 = frame (4k)
frame_vm_group_bin_13569 = frame (4k)
frame_vm_group_bin_1357 = frame (4k)
frame_vm_group_bin_13570 = frame (4k)
frame_vm_group_bin_13571 = frame (4k)
frame_vm_group_bin_13572 = frame (4k)
frame_vm_group_bin_13573 = frame (4k)
frame_vm_group_bin_13574 = frame (4k)
frame_vm_group_bin_13575 = frame (4k)
frame_vm_group_bin_13576 = frame (4k)
frame_vm_group_bin_13577 = frame (4k)
frame_vm_group_bin_13578 = frame (4k)
frame_vm_group_bin_13579 = frame (4k)
frame_vm_group_bin_1358 = frame (4k)
frame_vm_group_bin_13580 = frame (4k)
frame_vm_group_bin_13581 = frame (4k)
frame_vm_group_bin_13582 = frame (4k)
frame_vm_group_bin_13583 = frame (4k)
frame_vm_group_bin_13584 = frame (4k)
frame_vm_group_bin_13585 = frame (4k)
frame_vm_group_bin_13586 = frame (4k)
frame_vm_group_bin_13587 = frame (4k)
frame_vm_group_bin_13588 = frame (4k)
frame_vm_group_bin_13589 = frame (4k)
frame_vm_group_bin_1359 = frame (4k)
frame_vm_group_bin_13590 = frame (4k)
frame_vm_group_bin_13591 = frame (4k)
frame_vm_group_bin_13592 = frame (4k)
frame_vm_group_bin_13593 = frame (4k)
frame_vm_group_bin_13594 = frame (4k)
frame_vm_group_bin_13595 = frame (4k)
frame_vm_group_bin_13596 = frame (4k)
frame_vm_group_bin_13597 = frame (4k)
frame_vm_group_bin_13598 = frame (4k)
frame_vm_group_bin_13599 = frame (4k)
frame_vm_group_bin_1360 = frame (4k)
frame_vm_group_bin_13600 = frame (4k)
frame_vm_group_bin_13601 = frame (4k)
frame_vm_group_bin_13602 = frame (4k)
frame_vm_group_bin_13603 = frame (4k)
frame_vm_group_bin_13604 = frame (4k)
frame_vm_group_bin_13605 = frame (4k)
frame_vm_group_bin_13606 = frame (4k)
frame_vm_group_bin_13607 = frame (4k)
frame_vm_group_bin_13608 = frame (4k)
frame_vm_group_bin_13609 = frame (4k)
frame_vm_group_bin_1361 = frame (4k)
frame_vm_group_bin_13610 = frame (4k)
frame_vm_group_bin_13611 = frame (4k)
frame_vm_group_bin_13612 = frame (4k)
frame_vm_group_bin_13613 = frame (4k)
frame_vm_group_bin_13614 = frame (4k)
frame_vm_group_bin_13615 = frame (4k)
frame_vm_group_bin_13616 = frame (4k)
frame_vm_group_bin_13617 = frame (4k)
frame_vm_group_bin_13618 = frame (4k)
frame_vm_group_bin_13619 = frame (4k)
frame_vm_group_bin_1362 = frame (4k)
frame_vm_group_bin_13620 = frame (4k)
frame_vm_group_bin_13621 = frame (4k)
frame_vm_group_bin_13622 = frame (4k)
frame_vm_group_bin_13623 = frame (4k)
frame_vm_group_bin_13624 = frame (4k)
frame_vm_group_bin_13625 = frame (4k)
frame_vm_group_bin_13626 = frame (4k)
frame_vm_group_bin_13627 = frame (4k)
frame_vm_group_bin_13628 = frame (4k)
frame_vm_group_bin_13629 = frame (4k)
frame_vm_group_bin_1363 = frame (4k)
frame_vm_group_bin_13630 = frame (4k)
frame_vm_group_bin_13631 = frame (4k)
frame_vm_group_bin_13632 = frame (4k)
frame_vm_group_bin_13633 = frame (4k)
frame_vm_group_bin_13634 = frame (4k)
frame_vm_group_bin_13635 = frame (4k)
frame_vm_group_bin_13636 = frame (4k)
frame_vm_group_bin_13637 = frame (4k)
frame_vm_group_bin_13638 = frame (4k)
frame_vm_group_bin_13639 = frame (4k)
frame_vm_group_bin_1364 = frame (4k)
frame_vm_group_bin_13640 = frame (4k)
frame_vm_group_bin_13641 = frame (4k)
frame_vm_group_bin_13642 = frame (4k)
frame_vm_group_bin_13643 = frame (4k)
frame_vm_group_bin_13644 = frame (4k)
frame_vm_group_bin_13645 = frame (4k)
frame_vm_group_bin_13646 = frame (4k)
frame_vm_group_bin_13647 = frame (4k)
frame_vm_group_bin_13648 = frame (4k)
frame_vm_group_bin_13649 = frame (4k)
frame_vm_group_bin_1365 = frame (4k)
frame_vm_group_bin_13650 = frame (4k)
frame_vm_group_bin_13651 = frame (4k)
frame_vm_group_bin_13652 = frame (4k)
frame_vm_group_bin_13653 = frame (4k)
frame_vm_group_bin_13654 = frame (4k)
frame_vm_group_bin_13655 = frame (4k)
frame_vm_group_bin_13656 = frame (4k)
frame_vm_group_bin_13657 = frame (4k)
frame_vm_group_bin_13658 = frame (4k)
frame_vm_group_bin_13659 = frame (4k)
frame_vm_group_bin_1366 = frame (4k)
frame_vm_group_bin_13660 = frame (4k)
frame_vm_group_bin_13661 = frame (4k)
frame_vm_group_bin_13662 = frame (4k)
frame_vm_group_bin_13663 = frame (4k)
frame_vm_group_bin_13664 = frame (4k)
frame_vm_group_bin_13665 = frame (4k)
frame_vm_group_bin_13666 = frame (4k)
frame_vm_group_bin_13667 = frame (4k)
frame_vm_group_bin_13668 = frame (4k)
frame_vm_group_bin_13669 = frame (4k)
frame_vm_group_bin_1367 = frame (4k)
frame_vm_group_bin_13670 = frame (4k)
frame_vm_group_bin_13671 = frame (4k)
frame_vm_group_bin_13672 = frame (4k)
frame_vm_group_bin_13673 = frame (4k)
frame_vm_group_bin_13674 = frame (4k)
frame_vm_group_bin_13675 = frame (4k)
frame_vm_group_bin_13676 = frame (4k)
frame_vm_group_bin_13677 = frame (4k)
frame_vm_group_bin_13678 = frame (4k)
frame_vm_group_bin_13679 = frame (4k)
frame_vm_group_bin_1368 = frame (4k)
frame_vm_group_bin_13680 = frame (4k)
frame_vm_group_bin_13681 = frame (4k)
frame_vm_group_bin_13682 = frame (4k)
frame_vm_group_bin_13683 = frame (4k)
frame_vm_group_bin_13684 = frame (4k)
frame_vm_group_bin_13685 = frame (4k)
frame_vm_group_bin_13686 = frame (4k)
frame_vm_group_bin_13687 = frame (4k)
frame_vm_group_bin_13688 = frame (4k)
frame_vm_group_bin_13689 = frame (4k)
frame_vm_group_bin_1369 = frame (4k)
frame_vm_group_bin_13690 = frame (4k)
frame_vm_group_bin_13691 = frame (4k)
frame_vm_group_bin_13692 = frame (4k)
frame_vm_group_bin_13693 = frame (4k)
frame_vm_group_bin_13694 = frame (4k)
frame_vm_group_bin_13695 = frame (4k)
frame_vm_group_bin_13696 = frame (4k)
frame_vm_group_bin_13697 = frame (4k)
frame_vm_group_bin_13698 = frame (4k)
frame_vm_group_bin_13699 = frame (4k)
frame_vm_group_bin_1370 = frame (4k)
frame_vm_group_bin_13700 = frame (4k)
frame_vm_group_bin_13701 = frame (4k)
frame_vm_group_bin_13702 = frame (4k)
frame_vm_group_bin_13703 = frame (4k)
frame_vm_group_bin_13704 = frame (4k)
frame_vm_group_bin_13705 = frame (4k)
frame_vm_group_bin_13706 = frame (4k)
frame_vm_group_bin_13707 = frame (4k)
frame_vm_group_bin_13708 = frame (4k)
frame_vm_group_bin_13709 = frame (4k)
frame_vm_group_bin_1371 = frame (4k)
frame_vm_group_bin_13710 = frame (4k)
frame_vm_group_bin_13711 = frame (4k)
frame_vm_group_bin_13712 = frame (4k)
frame_vm_group_bin_13713 = frame (4k)
frame_vm_group_bin_13714 = frame (4k)
frame_vm_group_bin_13715 = frame (4k)
frame_vm_group_bin_13716 = frame (4k)
frame_vm_group_bin_13717 = frame (4k)
frame_vm_group_bin_13718 = frame (4k)
frame_vm_group_bin_13719 = frame (4k)
frame_vm_group_bin_1372 = frame (4k)
frame_vm_group_bin_13720 = frame (4k)
frame_vm_group_bin_13721 = frame (4k)
frame_vm_group_bin_13722 = frame (4k)
frame_vm_group_bin_13723 = frame (4k)
frame_vm_group_bin_13724 = frame (4k)
frame_vm_group_bin_13725 = frame (4k)
frame_vm_group_bin_13726 = frame (4k)
frame_vm_group_bin_13727 = frame (4k)
frame_vm_group_bin_13728 = frame (4k)
frame_vm_group_bin_13729 = frame (4k)
frame_vm_group_bin_1373 = frame (4k)
frame_vm_group_bin_13730 = frame (4k)
frame_vm_group_bin_13731 = frame (4k)
frame_vm_group_bin_13732 = frame (4k)
frame_vm_group_bin_13733 = frame (4k)
frame_vm_group_bin_13734 = frame (4k)
frame_vm_group_bin_13735 = frame (4k)
frame_vm_group_bin_13736 = frame (4k)
frame_vm_group_bin_13737 = frame (4k)
frame_vm_group_bin_13738 = frame (4k)
frame_vm_group_bin_13739 = frame (4k)
frame_vm_group_bin_1374 = frame (4k)
frame_vm_group_bin_13740 = frame (4k)
frame_vm_group_bin_13741 = frame (4k)
frame_vm_group_bin_13742 = frame (4k)
frame_vm_group_bin_13743 = frame (4k)
frame_vm_group_bin_13744 = frame (4k)
frame_vm_group_bin_13745 = frame (4k)
frame_vm_group_bin_13746 = frame (4k)
frame_vm_group_bin_13747 = frame (4k)
frame_vm_group_bin_13748 = frame (4k)
frame_vm_group_bin_13749 = frame (4k)
frame_vm_group_bin_1375 = frame (4k)
frame_vm_group_bin_13750 = frame (4k)
frame_vm_group_bin_13751 = frame (4k)
frame_vm_group_bin_13752 = frame (4k)
frame_vm_group_bin_13753 = frame (4k)
frame_vm_group_bin_13754 = frame (4k)
frame_vm_group_bin_13755 = frame (4k)
frame_vm_group_bin_13756 = frame (4k)
frame_vm_group_bin_13757 = frame (4k)
frame_vm_group_bin_13758 = frame (4k)
frame_vm_group_bin_13759 = frame (4k)
frame_vm_group_bin_1376 = frame (4k)
frame_vm_group_bin_13760 = frame (4k)
frame_vm_group_bin_13761 = frame (4k)
frame_vm_group_bin_13762 = frame (4k)
frame_vm_group_bin_13763 = frame (4k)
frame_vm_group_bin_13764 = frame (4k)
frame_vm_group_bin_13765 = frame (4k)
frame_vm_group_bin_13766 = frame (4k)
frame_vm_group_bin_13767 = frame (4k)
frame_vm_group_bin_13768 = frame (4k)
frame_vm_group_bin_13769 = frame (4k)
frame_vm_group_bin_1377 = frame (4k)
frame_vm_group_bin_13770 = frame (4k)
frame_vm_group_bin_13771 = frame (4k)
frame_vm_group_bin_13772 = frame (4k)
frame_vm_group_bin_13773 = frame (4k)
frame_vm_group_bin_13774 = frame (4k)
frame_vm_group_bin_13775 = frame (4k)
frame_vm_group_bin_13776 = frame (4k)
frame_vm_group_bin_13777 = frame (4k)
frame_vm_group_bin_13778 = frame (4k)
frame_vm_group_bin_13779 = frame (4k)
frame_vm_group_bin_1378 = frame (4k)
frame_vm_group_bin_13780 = frame (4k)
frame_vm_group_bin_13781 = frame (4k)
frame_vm_group_bin_13782 = frame (4k)
frame_vm_group_bin_13783 = frame (4k)
frame_vm_group_bin_13784 = frame (4k)
frame_vm_group_bin_13785 = frame (4k)
frame_vm_group_bin_13786 = frame (4k)
frame_vm_group_bin_13787 = frame (4k)
frame_vm_group_bin_13788 = frame (4k)
frame_vm_group_bin_13789 = frame (4k)
frame_vm_group_bin_1379 = frame (4k)
frame_vm_group_bin_13790 = frame (4k)
frame_vm_group_bin_13791 = frame (4k)
frame_vm_group_bin_13792 = frame (4k)
frame_vm_group_bin_13793 = frame (4k)
frame_vm_group_bin_13794 = frame (4k)
frame_vm_group_bin_13795 = frame (4k)
frame_vm_group_bin_13796 = frame (4k)
frame_vm_group_bin_13797 = frame (4k)
frame_vm_group_bin_13798 = frame (4k)
frame_vm_group_bin_13799 = frame (4k)
frame_vm_group_bin_1380 = frame (4k)
frame_vm_group_bin_13800 = frame (4k)
frame_vm_group_bin_13801 = frame (4k)
frame_vm_group_bin_13802 = frame (4k)
frame_vm_group_bin_13803 = frame (4k)
frame_vm_group_bin_13804 = frame (4k)
frame_vm_group_bin_13805 = frame (4k)
frame_vm_group_bin_13806 = frame (4k)
frame_vm_group_bin_13807 = frame (4k)
frame_vm_group_bin_13808 = frame (4k)
frame_vm_group_bin_13809 = frame (4k)
frame_vm_group_bin_1381 = frame (4k)
frame_vm_group_bin_13810 = frame (4k)
frame_vm_group_bin_13811 = frame (4k)
frame_vm_group_bin_13812 = frame (4k)
frame_vm_group_bin_13813 = frame (4k)
frame_vm_group_bin_13814 = frame (4k)
frame_vm_group_bin_13815 = frame (4k)
frame_vm_group_bin_13816 = frame (4k)
frame_vm_group_bin_13817 = frame (4k)
frame_vm_group_bin_13818 = frame (4k)
frame_vm_group_bin_13819 = frame (4k)
frame_vm_group_bin_1382 = frame (4k)
frame_vm_group_bin_13820 = frame (4k)
frame_vm_group_bin_13821 = frame (4k)
frame_vm_group_bin_13822 = frame (4k)
frame_vm_group_bin_13823 = frame (4k)
frame_vm_group_bin_13824 = frame (4k)
frame_vm_group_bin_13825 = frame (4k)
frame_vm_group_bin_13826 = frame (4k)
frame_vm_group_bin_13827 = frame (4k)
frame_vm_group_bin_13828 = frame (4k)
frame_vm_group_bin_13829 = frame (4k)
frame_vm_group_bin_1383 = frame (4k)
frame_vm_group_bin_13830 = frame (4k)
frame_vm_group_bin_13831 = frame (4k)
frame_vm_group_bin_13832 = frame (4k)
frame_vm_group_bin_13833 = frame (4k)
frame_vm_group_bin_13834 = frame (4k)
frame_vm_group_bin_13835 = frame (4k)
frame_vm_group_bin_13836 = frame (4k)
frame_vm_group_bin_13837 = frame (4k)
frame_vm_group_bin_13838 = frame (4k)
frame_vm_group_bin_13839 = frame (4k)
frame_vm_group_bin_1384 = frame (4k)
frame_vm_group_bin_13840 = frame (4k)
frame_vm_group_bin_13841 = frame (4k)
frame_vm_group_bin_13842 = frame (4k)
frame_vm_group_bin_13843 = frame (4k)
frame_vm_group_bin_13844 = frame (4k)
frame_vm_group_bin_13845 = frame (4k)
frame_vm_group_bin_13846 = frame (4k)
frame_vm_group_bin_13847 = frame (4k)
frame_vm_group_bin_13848 = frame (4k)
frame_vm_group_bin_13849 = frame (4k)
frame_vm_group_bin_1385 = frame (4k)
frame_vm_group_bin_13850 = frame (4k)
frame_vm_group_bin_13851 = frame (4k)
frame_vm_group_bin_13852 = frame (4k)
frame_vm_group_bin_13853 = frame (4k)
frame_vm_group_bin_13854 = frame (4k)
frame_vm_group_bin_13855 = frame (4k)
frame_vm_group_bin_13856 = frame (4k)
frame_vm_group_bin_13857 = frame (4k)
frame_vm_group_bin_13858 = frame (4k)
frame_vm_group_bin_13859 = frame (4k)
frame_vm_group_bin_1386 = frame (4k)
frame_vm_group_bin_13860 = frame (4k)
frame_vm_group_bin_13861 = frame (4k)
frame_vm_group_bin_13862 = frame (4k)
frame_vm_group_bin_13863 = frame (4k)
frame_vm_group_bin_13864 = frame (4k)
frame_vm_group_bin_13865 = frame (4k)
frame_vm_group_bin_13866 = frame (4k)
frame_vm_group_bin_13867 = frame (4k)
frame_vm_group_bin_13868 = frame (4k)
frame_vm_group_bin_13869 = frame (4k)
frame_vm_group_bin_1387 = frame (4k)
frame_vm_group_bin_13870 = frame (4k)
frame_vm_group_bin_13871 = frame (4k)
frame_vm_group_bin_13872 = frame (4k)
frame_vm_group_bin_13873 = frame (4k)
frame_vm_group_bin_13874 = frame (4k)
frame_vm_group_bin_13875 = frame (4k)
frame_vm_group_bin_13876 = frame (4k)
frame_vm_group_bin_13877 = frame (4k)
frame_vm_group_bin_13878 = frame (4k)
frame_vm_group_bin_13879 = frame (4k)
frame_vm_group_bin_1388 = frame (4k)
frame_vm_group_bin_13880 = frame (4k)
frame_vm_group_bin_13881 = frame (4k)
frame_vm_group_bin_13882 = frame (4k)
frame_vm_group_bin_13883 = frame (4k)
frame_vm_group_bin_13884 = frame (4k)
frame_vm_group_bin_13885 = frame (4k)
frame_vm_group_bin_13886 = frame (4k)
frame_vm_group_bin_13887 = frame (4k)
frame_vm_group_bin_13888 = frame (4k)
frame_vm_group_bin_13889 = frame (4k)
frame_vm_group_bin_1389 = frame (4k)
frame_vm_group_bin_13890 = frame (4k)
frame_vm_group_bin_13891 = frame (4k)
frame_vm_group_bin_13892 = frame (4k)
frame_vm_group_bin_13893 = frame (4k)
frame_vm_group_bin_13894 = frame (4k)
frame_vm_group_bin_13895 = frame (4k)
frame_vm_group_bin_13896 = frame (4k)
frame_vm_group_bin_13897 = frame (4k)
frame_vm_group_bin_13898 = frame (4k)
frame_vm_group_bin_13899 = frame (4k)
frame_vm_group_bin_1390 = frame (4k)
frame_vm_group_bin_13900 = frame (4k)
frame_vm_group_bin_13901 = frame (4k)
frame_vm_group_bin_13902 = frame (4k)
frame_vm_group_bin_13903 = frame (4k)
frame_vm_group_bin_13904 = frame (4k)
frame_vm_group_bin_13905 = frame (4k)
frame_vm_group_bin_13906 = frame (4k)
frame_vm_group_bin_13907 = frame (4k)
frame_vm_group_bin_13908 = frame (4k)
frame_vm_group_bin_13909 = frame (4k)
frame_vm_group_bin_1391 = frame (4k)
frame_vm_group_bin_13910 = frame (4k)
frame_vm_group_bin_13911 = frame (4k)
frame_vm_group_bin_13912 = frame (4k)
frame_vm_group_bin_13913 = frame (4k)
frame_vm_group_bin_13914 = frame (4k)
frame_vm_group_bin_13915 = frame (4k)
frame_vm_group_bin_13916 = frame (4k)
frame_vm_group_bin_13917 = frame (4k)
frame_vm_group_bin_13918 = frame (4k)
frame_vm_group_bin_13919 = frame (4k)
frame_vm_group_bin_1392 = frame (4k)
frame_vm_group_bin_13920 = frame (4k)
frame_vm_group_bin_13921 = frame (4k)
frame_vm_group_bin_13922 = frame (4k)
frame_vm_group_bin_13923 = frame (4k)
frame_vm_group_bin_13924 = frame (4k)
frame_vm_group_bin_13925 = frame (4k)
frame_vm_group_bin_13926 = frame (4k)
frame_vm_group_bin_13927 = frame (4k)
frame_vm_group_bin_13928 = frame (4k)
frame_vm_group_bin_13929 = frame (4k)
frame_vm_group_bin_1393 = frame (4k)
frame_vm_group_bin_13930 = frame (4k)
frame_vm_group_bin_13931 = frame (4k)
frame_vm_group_bin_13932 = frame (4k)
frame_vm_group_bin_13933 = frame (4k)
frame_vm_group_bin_13934 = frame (4k)
frame_vm_group_bin_13935 = frame (4k)
frame_vm_group_bin_13936 = frame (4k)
frame_vm_group_bin_13937 = frame (4k)
frame_vm_group_bin_13938 = frame (4k)
frame_vm_group_bin_13939 = frame (4k)
frame_vm_group_bin_1394 = frame (4k)
frame_vm_group_bin_13940 = frame (4k)
frame_vm_group_bin_13941 = frame (4k)
frame_vm_group_bin_13942 = frame (4k)
frame_vm_group_bin_13943 = frame (4k)
frame_vm_group_bin_13944 = frame (4k)
frame_vm_group_bin_13945 = frame (4k)
frame_vm_group_bin_13946 = frame (4k)
frame_vm_group_bin_13947 = frame (4k)
frame_vm_group_bin_13948 = frame (4k)
frame_vm_group_bin_13949 = frame (4k)
frame_vm_group_bin_1395 = frame (4k)
frame_vm_group_bin_13950 = frame (4k)
frame_vm_group_bin_13951 = frame (4k)
frame_vm_group_bin_13952 = frame (4k)
frame_vm_group_bin_13953 = frame (4k)
frame_vm_group_bin_13954 = frame (4k)
frame_vm_group_bin_13955 = frame (4k)
frame_vm_group_bin_13956 = frame (4k)
frame_vm_group_bin_13957 = frame (4k)
frame_vm_group_bin_13958 = frame (4k)
frame_vm_group_bin_13959 = frame (4k)
frame_vm_group_bin_1396 = frame (4k)
frame_vm_group_bin_13960 = frame (4k)
frame_vm_group_bin_13961 = frame (4k)
frame_vm_group_bin_13962 = frame (4k)
frame_vm_group_bin_13963 = frame (4k)
frame_vm_group_bin_13964 = frame (4k)
frame_vm_group_bin_13965 = frame (4k)
frame_vm_group_bin_13966 = frame (4k)
frame_vm_group_bin_13967 = frame (4k)
frame_vm_group_bin_13968 = frame (4k)
frame_vm_group_bin_13969 = frame (4k)
frame_vm_group_bin_1397 = frame (4k)
frame_vm_group_bin_13970 = frame (4k)
frame_vm_group_bin_13971 = frame (4k)
frame_vm_group_bin_13972 = frame (4k)
frame_vm_group_bin_13973 = frame (4k)
frame_vm_group_bin_13974 = frame (4k)
frame_vm_group_bin_13975 = frame (4k)
frame_vm_group_bin_13976 = frame (4k)
frame_vm_group_bin_13977 = frame (4k)
frame_vm_group_bin_13978 = frame (4k)
frame_vm_group_bin_13979 = frame (4k)
frame_vm_group_bin_1398 = frame (4k)
frame_vm_group_bin_13980 = frame (4k)
frame_vm_group_bin_13981 = frame (4k)
frame_vm_group_bin_13982 = frame (4k)
frame_vm_group_bin_13983 = frame (4k)
frame_vm_group_bin_13984 = frame (4k)
frame_vm_group_bin_13985 = frame (4k)
frame_vm_group_bin_13986 = frame (4k)
frame_vm_group_bin_13987 = frame (4k)
frame_vm_group_bin_13988 = frame (4k)
frame_vm_group_bin_13989 = frame (4k)
frame_vm_group_bin_1399 = frame (4k)
frame_vm_group_bin_13990 = frame (4k)
frame_vm_group_bin_13991 = frame (4k)
frame_vm_group_bin_13992 = frame (4k)
frame_vm_group_bin_13993 = frame (4k)
frame_vm_group_bin_13994 = frame (4k)
frame_vm_group_bin_13995 = frame (4k)
frame_vm_group_bin_13996 = frame (4k)
frame_vm_group_bin_13997 = frame (4k)
frame_vm_group_bin_13998 = frame (4k)
frame_vm_group_bin_13999 = frame (4k)
frame_vm_group_bin_1400 = frame (4k)
frame_vm_group_bin_14000 = frame (4k)
frame_vm_group_bin_14001 = frame (4k)
frame_vm_group_bin_14002 = frame (4k)
frame_vm_group_bin_14003 = frame (4k)
frame_vm_group_bin_14004 = frame (4k)
frame_vm_group_bin_14005 = frame (4k)
frame_vm_group_bin_14006 = frame (4k)
frame_vm_group_bin_14007 = frame (4k)
frame_vm_group_bin_14008 = frame (4k)
frame_vm_group_bin_14009 = frame (4k)
frame_vm_group_bin_1401 = frame (4k)
frame_vm_group_bin_14010 = frame (4k)
frame_vm_group_bin_14011 = frame (4k)
frame_vm_group_bin_14012 = frame (4k)
frame_vm_group_bin_14013 = frame (4k)
frame_vm_group_bin_14014 = frame (4k)
frame_vm_group_bin_14015 = frame (4k)
frame_vm_group_bin_14016 = frame (4k)
frame_vm_group_bin_14017 = frame (4k)
frame_vm_group_bin_14018 = frame (4k)
frame_vm_group_bin_14019 = frame (4k)
frame_vm_group_bin_1402 = frame (4k)
frame_vm_group_bin_14020 = frame (4k)
frame_vm_group_bin_14021 = frame (4k)
frame_vm_group_bin_14022 = frame (4k)
frame_vm_group_bin_14023 = frame (4k)
frame_vm_group_bin_14024 = frame (4k)
frame_vm_group_bin_14025 = frame (4k)
frame_vm_group_bin_14026 = frame (4k)
frame_vm_group_bin_14027 = frame (4k)
frame_vm_group_bin_14028 = frame (4k)
frame_vm_group_bin_14029 = frame (4k)
frame_vm_group_bin_1403 = frame (4k)
frame_vm_group_bin_14030 = frame (4k)
frame_vm_group_bin_14031 = frame (4k)
frame_vm_group_bin_14032 = frame (4k)
frame_vm_group_bin_14033 = frame (4k)
frame_vm_group_bin_14034 = frame (4k)
frame_vm_group_bin_14035 = frame (4k)
frame_vm_group_bin_14036 = frame (4k)
frame_vm_group_bin_14037 = frame (4k)
frame_vm_group_bin_14038 = frame (4k)
frame_vm_group_bin_14039 = frame (4k)
frame_vm_group_bin_1404 = frame (4k)
frame_vm_group_bin_14040 = frame (4k)
frame_vm_group_bin_14041 = frame (4k)
frame_vm_group_bin_14042 = frame (4k)
frame_vm_group_bin_14043 = frame (4k)
frame_vm_group_bin_14044 = frame (4k)
frame_vm_group_bin_14045 = frame (4k)
frame_vm_group_bin_14046 = frame (4k)
frame_vm_group_bin_14047 = frame (4k)
frame_vm_group_bin_14048 = frame (4k)
frame_vm_group_bin_14049 = frame (4k)
frame_vm_group_bin_1405 = frame (4k)
frame_vm_group_bin_14050 = frame (4k)
frame_vm_group_bin_14051 = frame (4k)
frame_vm_group_bin_14052 = frame (4k)
frame_vm_group_bin_14053 = frame (4k)
frame_vm_group_bin_14054 = frame (4k)
frame_vm_group_bin_14055 = frame (4k)
frame_vm_group_bin_14056 = frame (4k)
frame_vm_group_bin_14057 = frame (4k)
frame_vm_group_bin_14058 = frame (4k)
frame_vm_group_bin_14059 = frame (4k)
frame_vm_group_bin_1406 = frame (4k)
frame_vm_group_bin_14060 = frame (4k)
frame_vm_group_bin_14061 = frame (4k)
frame_vm_group_bin_14062 = frame (4k)
frame_vm_group_bin_14063 = frame (4k)
frame_vm_group_bin_14064 = frame (4k)
frame_vm_group_bin_14065 = frame (4k)
frame_vm_group_bin_14066 = frame (4k)
frame_vm_group_bin_14067 = frame (4k)
frame_vm_group_bin_14068 = frame (4k)
frame_vm_group_bin_14069 = frame (4k)
frame_vm_group_bin_1407 = frame (4k)
frame_vm_group_bin_14070 = frame (4k)
frame_vm_group_bin_14071 = frame (4k)
frame_vm_group_bin_14072 = frame (4k)
frame_vm_group_bin_14073 = frame (4k)
frame_vm_group_bin_14074 = frame (4k)
frame_vm_group_bin_14075 = frame (4k)
frame_vm_group_bin_14076 = frame (4k)
frame_vm_group_bin_14077 = frame (4k)
frame_vm_group_bin_14078 = frame (4k)
frame_vm_group_bin_14079 = frame (4k)
frame_vm_group_bin_1408 = frame (4k)
frame_vm_group_bin_14080 = frame (4k)
frame_vm_group_bin_14081 = frame (4k)
frame_vm_group_bin_14082 = frame (4k)
frame_vm_group_bin_14083 = frame (4k)
frame_vm_group_bin_14084 = frame (4k)
frame_vm_group_bin_14085 = frame (4k)
frame_vm_group_bin_14086 = frame (4k)
frame_vm_group_bin_14087 = frame (4k)
frame_vm_group_bin_14088 = frame (4k)
frame_vm_group_bin_14089 = frame (4k)
frame_vm_group_bin_1409 = frame (4k)
frame_vm_group_bin_14090 = frame (4k)
frame_vm_group_bin_14091 = frame (4k)
frame_vm_group_bin_14092 = frame (4k)
frame_vm_group_bin_14093 = frame (4k)
frame_vm_group_bin_14094 = frame (4k)
frame_vm_group_bin_14095 = frame (4k)
frame_vm_group_bin_14096 = frame (4k)
frame_vm_group_bin_14097 = frame (4k)
frame_vm_group_bin_14098 = frame (4k)
frame_vm_group_bin_14099 = frame (4k)
frame_vm_group_bin_1410 = frame (4k)
frame_vm_group_bin_14100 = frame (4k)
frame_vm_group_bin_14101 = frame (4k)
frame_vm_group_bin_14102 = frame (4k)
frame_vm_group_bin_14103 = frame (4k)
frame_vm_group_bin_14104 = frame (4k)
frame_vm_group_bin_14105 = frame (4k)
frame_vm_group_bin_14106 = frame (4k)
frame_vm_group_bin_14107 = frame (4k)
frame_vm_group_bin_14108 = frame (4k)
frame_vm_group_bin_14109 = frame (4k)
frame_vm_group_bin_1411 = frame (4k)
frame_vm_group_bin_14110 = frame (4k)
frame_vm_group_bin_14111 = frame (4k)
frame_vm_group_bin_14112 = frame (4k)
frame_vm_group_bin_14113 = frame (4k)
frame_vm_group_bin_14114 = frame (4k)
frame_vm_group_bin_14115 = frame (4k)
frame_vm_group_bin_14116 = frame (4k)
frame_vm_group_bin_14117 = frame (4k)
frame_vm_group_bin_14118 = frame (4k)
frame_vm_group_bin_14119 = frame (4k)
frame_vm_group_bin_1412 = frame (4k)
frame_vm_group_bin_14120 = frame (4k)
frame_vm_group_bin_14121 = frame (4k)
frame_vm_group_bin_14122 = frame (4k)
frame_vm_group_bin_14123 = frame (4k)
frame_vm_group_bin_14124 = frame (4k)
frame_vm_group_bin_14125 = frame (4k)
frame_vm_group_bin_14126 = frame (4k)
frame_vm_group_bin_14127 = frame (4k)
frame_vm_group_bin_14128 = frame (4k)
frame_vm_group_bin_14129 = frame (4k)
frame_vm_group_bin_1413 = frame (4k)
frame_vm_group_bin_14130 = frame (4k)
frame_vm_group_bin_14131 = frame (4k)
frame_vm_group_bin_14132 = frame (4k)
frame_vm_group_bin_14133 = frame (4k)
frame_vm_group_bin_14134 = frame (4k)
frame_vm_group_bin_14135 = frame (4k)
frame_vm_group_bin_14136 = frame (4k)
frame_vm_group_bin_14137 = frame (4k)
frame_vm_group_bin_14138 = frame (4k)
frame_vm_group_bin_14139 = frame (4k)
frame_vm_group_bin_1414 = frame (4k)
frame_vm_group_bin_14140 = frame (4k)
frame_vm_group_bin_14141 = frame (4k)
frame_vm_group_bin_14142 = frame (4k)
frame_vm_group_bin_14143 = frame (4k)
frame_vm_group_bin_14144 = frame (4k)
frame_vm_group_bin_14145 = frame (4k)
frame_vm_group_bin_14146 = frame (4k)
frame_vm_group_bin_14147 = frame (4k)
frame_vm_group_bin_14148 = frame (4k)
frame_vm_group_bin_14149 = frame (4k)
frame_vm_group_bin_1415 = frame (4k)
frame_vm_group_bin_14150 = frame (4k)
frame_vm_group_bin_14151 = frame (4k)
frame_vm_group_bin_14152 = frame (4k)
frame_vm_group_bin_14153 = frame (4k)
frame_vm_group_bin_14154 = frame (4k)
frame_vm_group_bin_14155 = frame (4k)
frame_vm_group_bin_14156 = frame (4k)
frame_vm_group_bin_14157 = frame (4k)
frame_vm_group_bin_14158 = frame (4k)
frame_vm_group_bin_14159 = frame (4k)
frame_vm_group_bin_1416 = frame (4k)
frame_vm_group_bin_14160 = frame (4k)
frame_vm_group_bin_14161 = frame (4k)
frame_vm_group_bin_14162 = frame (4k)
frame_vm_group_bin_14163 = frame (4k)
frame_vm_group_bin_14164 = frame (4k)
frame_vm_group_bin_14165 = frame (4k)
frame_vm_group_bin_14166 = frame (4k)
frame_vm_group_bin_14167 = frame (4k)
frame_vm_group_bin_14168 = frame (4k)
frame_vm_group_bin_14169 = frame (4k)
frame_vm_group_bin_1417 = frame (4k)
frame_vm_group_bin_14170 = frame (4k)
frame_vm_group_bin_14171 = frame (4k)
frame_vm_group_bin_14172 = frame (4k)
frame_vm_group_bin_14173 = frame (4k)
frame_vm_group_bin_14174 = frame (4k)
frame_vm_group_bin_14175 = frame (4k)
frame_vm_group_bin_14176 = frame (4k)
frame_vm_group_bin_14177 = frame (4k)
frame_vm_group_bin_14178 = frame (4k)
frame_vm_group_bin_14179 = frame (4k)
frame_vm_group_bin_1418 = frame (4k)
frame_vm_group_bin_14180 = frame (4k)
frame_vm_group_bin_14182 = frame (4k)
frame_vm_group_bin_14183 = frame (4k)
frame_vm_group_bin_14184 = frame (4k)
frame_vm_group_bin_14185 = frame (4k)
frame_vm_group_bin_14186 = frame (4k)
frame_vm_group_bin_14187 = frame (4k)
frame_vm_group_bin_14188 = frame (4k)
frame_vm_group_bin_14189 = frame (4k)
frame_vm_group_bin_1419 = frame (4k)
frame_vm_group_bin_14190 = frame (4k)
frame_vm_group_bin_14191 = frame (4k)
frame_vm_group_bin_14192 = frame (4k)
frame_vm_group_bin_14193 = frame (4k)
frame_vm_group_bin_14194 = frame (4k)
frame_vm_group_bin_14195 = frame (4k)
frame_vm_group_bin_14196 = frame (4k)
frame_vm_group_bin_14197 = frame (4k)
frame_vm_group_bin_14198 = frame (4k)
frame_vm_group_bin_14199 = frame (4k)
frame_vm_group_bin_1420 = frame (4k)
frame_vm_group_bin_14200 = frame (4k)
frame_vm_group_bin_14201 = frame (4k)
frame_vm_group_bin_14202 = frame (4k)
frame_vm_group_bin_14203 = frame (4k)
frame_vm_group_bin_14204 = frame (4k)
frame_vm_group_bin_14205 = frame (4k)
frame_vm_group_bin_14206 = frame (4k)
frame_vm_group_bin_14207 = frame (4k)
frame_vm_group_bin_14208 = frame (4k)
frame_vm_group_bin_14209 = frame (4k)
frame_vm_group_bin_1421 = frame (4k)
frame_vm_group_bin_14210 = frame (4k)
frame_vm_group_bin_14211 = frame (4k)
frame_vm_group_bin_14212 = frame (4k)
frame_vm_group_bin_14213 = frame (4k)
frame_vm_group_bin_14214 = frame (4k)
frame_vm_group_bin_14215 = frame (4k)
frame_vm_group_bin_14216 = frame (4k)
frame_vm_group_bin_14217 = frame (4k)
frame_vm_group_bin_14218 = frame (4k)
frame_vm_group_bin_14219 = frame (4k)
frame_vm_group_bin_1422 = frame (4k)
frame_vm_group_bin_14220 = frame (4k)
frame_vm_group_bin_14221 = frame (4k)
frame_vm_group_bin_14222 = frame (4k)
frame_vm_group_bin_14223 = frame (4k)
frame_vm_group_bin_14224 = frame (4k)
frame_vm_group_bin_14225 = frame (4k)
frame_vm_group_bin_14226 = frame (4k)
frame_vm_group_bin_14227 = frame (4k)
frame_vm_group_bin_14228 = frame (4k)
frame_vm_group_bin_14229 = frame (4k)
frame_vm_group_bin_1423 = frame (4k)
frame_vm_group_bin_14230 = frame (4k)
frame_vm_group_bin_14231 = frame (4k)
frame_vm_group_bin_14232 = frame (4k)
frame_vm_group_bin_14233 = frame (4k)
frame_vm_group_bin_14234 = frame (4k)
frame_vm_group_bin_14235 = frame (4k)
frame_vm_group_bin_14236 = frame (4k)
frame_vm_group_bin_14237 = frame (4k)
frame_vm_group_bin_14238 = frame (4k)
frame_vm_group_bin_14239 = frame (4k)
frame_vm_group_bin_1424 = frame (4k)
frame_vm_group_bin_14240 = frame (4k)
frame_vm_group_bin_14241 = frame (4k)
frame_vm_group_bin_14242 = frame (4k)
frame_vm_group_bin_14243 = frame (4k)
frame_vm_group_bin_14244 = frame (4k)
frame_vm_group_bin_14245 = frame (4k)
frame_vm_group_bin_14246 = frame (4k)
frame_vm_group_bin_14247 = frame (4k)
frame_vm_group_bin_14248 = frame (4k)
frame_vm_group_bin_14249 = frame (4k)
frame_vm_group_bin_1425 = frame (4k)
frame_vm_group_bin_14250 = frame (4k)
frame_vm_group_bin_14251 = frame (4k)
frame_vm_group_bin_14252 = frame (4k)
frame_vm_group_bin_14253 = frame (4k)
frame_vm_group_bin_14254 = frame (4k)
frame_vm_group_bin_14255 = frame (4k)
frame_vm_group_bin_14256 = frame (4k)
frame_vm_group_bin_14257 = frame (4k)
frame_vm_group_bin_14258 = frame (4k)
frame_vm_group_bin_14259 = frame (4k)
frame_vm_group_bin_1426 = frame (4k)
frame_vm_group_bin_14260 = frame (4k)
frame_vm_group_bin_14261 = frame (4k)
frame_vm_group_bin_14262 = frame (4k)
frame_vm_group_bin_14263 = frame (4k)
frame_vm_group_bin_14264 = frame (4k)
frame_vm_group_bin_14265 = frame (4k)
frame_vm_group_bin_14266 = frame (4k)
frame_vm_group_bin_14267 = frame (4k)
frame_vm_group_bin_14268 = frame (4k)
frame_vm_group_bin_14269 = frame (4k)
frame_vm_group_bin_1427 = frame (4k)
frame_vm_group_bin_14270 = frame (4k)
frame_vm_group_bin_14271 = frame (4k)
frame_vm_group_bin_14272 = frame (4k)
frame_vm_group_bin_14273 = frame (4k)
frame_vm_group_bin_14274 = frame (4k)
frame_vm_group_bin_14275 = frame (4k)
frame_vm_group_bin_14276 = frame (4k)
frame_vm_group_bin_14277 = frame (4k)
frame_vm_group_bin_14278 = frame (4k)
frame_vm_group_bin_14279 = frame (4k)
frame_vm_group_bin_1428 = frame (4k)
frame_vm_group_bin_14280 = frame (4k)
frame_vm_group_bin_14281 = frame (4k)
frame_vm_group_bin_14282 = frame (4k)
frame_vm_group_bin_14283 = frame (4k)
frame_vm_group_bin_14284 = frame (4k)
frame_vm_group_bin_14285 = frame (4k)
frame_vm_group_bin_14286 = frame (4k)
frame_vm_group_bin_14287 = frame (4k)
frame_vm_group_bin_14288 = frame (4k)
frame_vm_group_bin_14289 = frame (4k)
frame_vm_group_bin_1429 = frame (4k)
frame_vm_group_bin_14290 = frame (4k)
frame_vm_group_bin_14291 = frame (4k)
frame_vm_group_bin_14292 = frame (4k)
frame_vm_group_bin_14293 = frame (4k)
frame_vm_group_bin_14294 = frame (4k)
frame_vm_group_bin_14295 = frame (4k)
frame_vm_group_bin_14296 = frame (4k)
frame_vm_group_bin_14297 = frame (4k)
frame_vm_group_bin_14298 = frame (4k)
frame_vm_group_bin_14299 = frame (4k)
frame_vm_group_bin_1430 = frame (4k)
frame_vm_group_bin_14300 = frame (4k)
frame_vm_group_bin_14301 = frame (4k)
frame_vm_group_bin_14302 = frame (4k)
frame_vm_group_bin_14303 = frame (4k)
frame_vm_group_bin_14304 = frame (4k)
frame_vm_group_bin_14305 = frame (4k)
frame_vm_group_bin_14306 = frame (4k)
frame_vm_group_bin_14307 = frame (4k)
frame_vm_group_bin_14308 = frame (4k)
frame_vm_group_bin_14309 = frame (4k)
frame_vm_group_bin_1431 = frame (4k)
frame_vm_group_bin_14310 = frame (4k)
frame_vm_group_bin_14311 = frame (4k)
frame_vm_group_bin_14312 = frame (4k)
frame_vm_group_bin_14313 = frame (4k)
frame_vm_group_bin_14314 = frame (4k)
frame_vm_group_bin_14315 = frame (4k)
frame_vm_group_bin_14316 = frame (4k)
frame_vm_group_bin_14317 = frame (4k)
frame_vm_group_bin_14318 = frame (4k)
frame_vm_group_bin_14319 = frame (4k)
frame_vm_group_bin_1432 = frame (4k)
frame_vm_group_bin_14320 = frame (4k)
frame_vm_group_bin_14321 = frame (4k)
frame_vm_group_bin_14322 = frame (4k)
frame_vm_group_bin_14323 = frame (4k)
frame_vm_group_bin_14324 = frame (4k)
frame_vm_group_bin_14325 = frame (4k)
frame_vm_group_bin_14326 = frame (4k)
frame_vm_group_bin_14327 = frame (4k)
frame_vm_group_bin_14328 = frame (4k)
frame_vm_group_bin_14329 = frame (4k)
frame_vm_group_bin_1433 = frame (4k)
frame_vm_group_bin_14330 = frame (4k)
frame_vm_group_bin_14331 = frame (4k)
frame_vm_group_bin_14332 = frame (4k)
frame_vm_group_bin_14333 = frame (4k)
frame_vm_group_bin_14334 = frame (4k)
frame_vm_group_bin_14335 = frame (4k)
frame_vm_group_bin_14336 = frame (4k)
frame_vm_group_bin_14337 = frame (4k)
frame_vm_group_bin_14338 = frame (4k)
frame_vm_group_bin_14339 = frame (4k)
frame_vm_group_bin_1434 = frame (4k)
frame_vm_group_bin_14340 = frame (4k)
frame_vm_group_bin_14341 = frame (4k)
frame_vm_group_bin_14342 = frame (4k)
frame_vm_group_bin_14343 = frame (4k)
frame_vm_group_bin_14344 = frame (4k)
frame_vm_group_bin_14345 = frame (4k)
frame_vm_group_bin_14346 = frame (4k)
frame_vm_group_bin_14347 = frame (4k)
frame_vm_group_bin_14348 = frame (4k)
frame_vm_group_bin_14349 = frame (4k)
frame_vm_group_bin_1435 = frame (4k)
frame_vm_group_bin_14350 = frame (4k)
frame_vm_group_bin_14351 = frame (4k)
frame_vm_group_bin_14352 = frame (4k)
frame_vm_group_bin_14353 = frame (4k)
frame_vm_group_bin_14354 = frame (4k)
frame_vm_group_bin_14355 = frame (4k)
frame_vm_group_bin_14356 = frame (4k)
frame_vm_group_bin_14357 = frame (4k)
frame_vm_group_bin_14358 = frame (4k)
frame_vm_group_bin_14359 = frame (4k)
frame_vm_group_bin_1436 = frame (4k)
frame_vm_group_bin_14360 = frame (4k)
frame_vm_group_bin_14361 = frame (4k)
frame_vm_group_bin_14362 = frame (4k)
frame_vm_group_bin_14363 = frame (4k)
frame_vm_group_bin_14364 = frame (4k)
frame_vm_group_bin_14365 = frame (4k)
frame_vm_group_bin_14366 = frame (4k)
frame_vm_group_bin_14367 = frame (4k)
frame_vm_group_bin_14368 = frame (4k)
frame_vm_group_bin_14369 = frame (4k)
frame_vm_group_bin_1437 = frame (4k)
frame_vm_group_bin_14370 = frame (4k)
frame_vm_group_bin_14371 = frame (4k)
frame_vm_group_bin_14372 = frame (4k)
frame_vm_group_bin_14373 = frame (4k)
frame_vm_group_bin_14374 = frame (4k)
frame_vm_group_bin_14375 = frame (4k)
frame_vm_group_bin_14376 = frame (4k)
frame_vm_group_bin_14377 = frame (4k)
frame_vm_group_bin_14378 = frame (4k)
frame_vm_group_bin_14379 = frame (4k)
frame_vm_group_bin_1438 = frame (4k)
frame_vm_group_bin_14380 = frame (4k)
frame_vm_group_bin_14381 = frame (4k)
frame_vm_group_bin_14382 = frame (4k)
frame_vm_group_bin_14383 = frame (4k)
frame_vm_group_bin_14384 = frame (4k)
frame_vm_group_bin_14385 = frame (4k)
frame_vm_group_bin_14386 = frame (4k)
frame_vm_group_bin_14387 = frame (4k)
frame_vm_group_bin_14388 = frame (4k)
frame_vm_group_bin_14389 = frame (4k)
frame_vm_group_bin_1439 = frame (4k)
frame_vm_group_bin_14390 = frame (4k)
frame_vm_group_bin_14391 = frame (4k)
frame_vm_group_bin_14392 = frame (4k)
frame_vm_group_bin_14393 = frame (4k)
frame_vm_group_bin_14394 = frame (4k)
frame_vm_group_bin_14395 = frame (4k)
frame_vm_group_bin_14396 = frame (4k)
frame_vm_group_bin_14397 = frame (4k)
frame_vm_group_bin_14398 = frame (4k)
frame_vm_group_bin_14399 = frame (4k)
frame_vm_group_bin_1440 = frame (4k)
frame_vm_group_bin_14400 = frame (4k)
frame_vm_group_bin_14401 = frame (4k)
frame_vm_group_bin_14402 = frame (4k)
frame_vm_group_bin_14403 = frame (4k)
frame_vm_group_bin_14404 = frame (4k)
frame_vm_group_bin_14405 = frame (4k)
frame_vm_group_bin_14406 = frame (4k)
frame_vm_group_bin_14407 = frame (4k)
frame_vm_group_bin_14408 = frame (4k)
frame_vm_group_bin_14409 = frame (4k)
frame_vm_group_bin_1441 = frame (4k)
frame_vm_group_bin_14410 = frame (4k)
frame_vm_group_bin_14411 = frame (4k)
frame_vm_group_bin_14412 = frame (4k)
frame_vm_group_bin_14413 = frame (4k)
frame_vm_group_bin_14414 = frame (4k)
frame_vm_group_bin_14415 = frame (4k)
frame_vm_group_bin_14416 = frame (4k)
frame_vm_group_bin_14417 = frame (4k)
frame_vm_group_bin_14418 = frame (4k)
frame_vm_group_bin_14419 = frame (4k)
frame_vm_group_bin_1442 = frame (4k)
frame_vm_group_bin_14420 = frame (4k)
frame_vm_group_bin_14421 = frame (4k)
frame_vm_group_bin_14422 = frame (4k)
frame_vm_group_bin_14423 = frame (4k)
frame_vm_group_bin_14424 = frame (4k)
frame_vm_group_bin_14425 = frame (4k)
frame_vm_group_bin_14426 = frame (4k)
frame_vm_group_bin_14427 = frame (4k)
frame_vm_group_bin_14428 = frame (4k)
frame_vm_group_bin_14429 = frame (4k)
frame_vm_group_bin_1443 = frame (4k)
frame_vm_group_bin_14430 = frame (4k)
frame_vm_group_bin_14431 = frame (4k)
frame_vm_group_bin_14432 = frame (4k)
frame_vm_group_bin_14433 = frame (4k)
frame_vm_group_bin_14434 = frame (4k)
frame_vm_group_bin_14435 = frame (4k)
frame_vm_group_bin_14436 = frame (4k)
frame_vm_group_bin_14437 = frame (4k)
frame_vm_group_bin_14438 = frame (4k)
frame_vm_group_bin_14439 = frame (4k)
frame_vm_group_bin_1444 = frame (4k)
frame_vm_group_bin_14440 = frame (4k)
frame_vm_group_bin_14441 = frame (4k)
frame_vm_group_bin_14442 = frame (4k)
frame_vm_group_bin_14443 = frame (4k)
frame_vm_group_bin_14444 = frame (4k)
frame_vm_group_bin_14445 = frame (4k)
frame_vm_group_bin_14446 = frame (4k)
frame_vm_group_bin_14447 = frame (4k)
frame_vm_group_bin_14448 = frame (4k)
frame_vm_group_bin_14449 = frame (4k)
frame_vm_group_bin_1445 = frame (4k)
frame_vm_group_bin_14450 = frame (4k)
frame_vm_group_bin_14451 = frame (4k)
frame_vm_group_bin_14452 = frame (4k)
frame_vm_group_bin_14453 = frame (4k)
frame_vm_group_bin_14454 = frame (4k)
frame_vm_group_bin_14455 = frame (4k)
frame_vm_group_bin_14456 = frame (4k)
frame_vm_group_bin_14457 = frame (4k)
frame_vm_group_bin_14458 = frame (4k)
frame_vm_group_bin_14459 = frame (4k)
frame_vm_group_bin_1446 = frame (4k)
frame_vm_group_bin_14460 = frame (4k)
frame_vm_group_bin_14461 = frame (4k)
frame_vm_group_bin_14462 = frame (4k)
frame_vm_group_bin_14463 = frame (4k)
frame_vm_group_bin_14464 = frame (4k)
frame_vm_group_bin_14465 = frame (4k)
frame_vm_group_bin_14466 = frame (4k)
frame_vm_group_bin_14467 = frame (4k)
frame_vm_group_bin_14468 = frame (4k)
frame_vm_group_bin_14469 = frame (4k)
frame_vm_group_bin_1447 = frame (4k)
frame_vm_group_bin_14470 = frame (4k)
frame_vm_group_bin_14471 = frame (4k)
frame_vm_group_bin_14472 = frame (4k)
frame_vm_group_bin_14473 = frame (4k)
frame_vm_group_bin_14474 = frame (4k)
frame_vm_group_bin_14475 = frame (4k)
frame_vm_group_bin_14476 = frame (4k)
frame_vm_group_bin_14477 = frame (4k)
frame_vm_group_bin_14478 = frame (4k)
frame_vm_group_bin_14479 = frame (4k)
frame_vm_group_bin_1448 = frame (4k)
frame_vm_group_bin_14480 = frame (4k)
frame_vm_group_bin_14481 = frame (4k)
frame_vm_group_bin_14482 = frame (4k)
frame_vm_group_bin_14483 = frame (4k)
frame_vm_group_bin_14484 = frame (4k)
frame_vm_group_bin_14485 = frame (4k)
frame_vm_group_bin_14486 = frame (4k)
frame_vm_group_bin_14487 = frame (4k)
frame_vm_group_bin_14488 = frame (4k)
frame_vm_group_bin_14489 = frame (4k)
frame_vm_group_bin_1449 = frame (4k)
frame_vm_group_bin_14490 = frame (4k)
frame_vm_group_bin_14491 = frame (4k)
frame_vm_group_bin_14492 = frame (4k)
frame_vm_group_bin_14493 = frame (4k)
frame_vm_group_bin_14494 = frame (4k)
frame_vm_group_bin_14495 = frame (4k)
frame_vm_group_bin_14496 = frame (4k)
frame_vm_group_bin_14497 = frame (4k)
frame_vm_group_bin_14498 = frame (4k)
frame_vm_group_bin_14499 = frame (4k)
frame_vm_group_bin_1450 = frame (4k)
frame_vm_group_bin_14500 = frame (4k)
frame_vm_group_bin_14501 = frame (4k)
frame_vm_group_bin_14502 = frame (4k)
frame_vm_group_bin_14503 = frame (4k)
frame_vm_group_bin_14504 = frame (4k)
frame_vm_group_bin_14505 = frame (4k)
frame_vm_group_bin_14506 = frame (4k)
frame_vm_group_bin_14507 = frame (4k)
frame_vm_group_bin_14508 = frame (4k)
frame_vm_group_bin_14509 = frame (4k)
frame_vm_group_bin_1451 = frame (4k)
frame_vm_group_bin_14510 = frame (4k)
frame_vm_group_bin_14511 = frame (4k)
frame_vm_group_bin_14512 = frame (4k)
frame_vm_group_bin_14513 = frame (4k)
frame_vm_group_bin_14514 = frame (4k)
frame_vm_group_bin_14515 = frame (4k)
frame_vm_group_bin_14516 = frame (4k)
frame_vm_group_bin_14517 = frame (4k)
frame_vm_group_bin_14518 = frame (4k)
frame_vm_group_bin_14519 = frame (4k)
frame_vm_group_bin_1452 = frame (4k)
frame_vm_group_bin_14520 = frame (4k)
frame_vm_group_bin_14521 = frame (4k)
frame_vm_group_bin_14522 = frame (4k)
frame_vm_group_bin_14523 = frame (4k)
frame_vm_group_bin_14524 = frame (4k)
frame_vm_group_bin_14525 = frame (4k)
frame_vm_group_bin_14526 = frame (4k)
frame_vm_group_bin_14527 = frame (4k)
frame_vm_group_bin_14528 = frame (4k)
frame_vm_group_bin_14529 = frame (4k)
frame_vm_group_bin_1453 = frame (4k)
frame_vm_group_bin_14530 = frame (4k)
frame_vm_group_bin_14531 = frame (4k)
frame_vm_group_bin_14532 = frame (4k)
frame_vm_group_bin_14533 = frame (4k)
frame_vm_group_bin_14534 = frame (4k)
frame_vm_group_bin_14535 = frame (4k)
frame_vm_group_bin_14536 = frame (4k)
frame_vm_group_bin_14537 = frame (4k)
frame_vm_group_bin_14538 = frame (4k)
frame_vm_group_bin_14539 = frame (4k)
frame_vm_group_bin_1454 = frame (4k)
frame_vm_group_bin_14540 = frame (4k)
frame_vm_group_bin_14541 = frame (4k)
frame_vm_group_bin_14542 = frame (4k)
frame_vm_group_bin_14543 = frame (4k)
frame_vm_group_bin_14544 = frame (4k)
frame_vm_group_bin_14545 = frame (4k)
frame_vm_group_bin_14546 = frame (4k)
frame_vm_group_bin_14547 = frame (4k)
frame_vm_group_bin_14548 = frame (4k)
frame_vm_group_bin_14549 = frame (4k)
frame_vm_group_bin_1455 = frame (4k)
frame_vm_group_bin_14550 = frame (4k)
frame_vm_group_bin_14551 = frame (4k)
frame_vm_group_bin_14552 = frame (4k)
frame_vm_group_bin_14553 = frame (4k)
frame_vm_group_bin_14554 = frame (4k)
frame_vm_group_bin_14555 = frame (4k)
frame_vm_group_bin_14556 = frame (4k)
frame_vm_group_bin_14557 = frame (4k)
frame_vm_group_bin_14558 = frame (4k)
frame_vm_group_bin_14559 = frame (4k)
frame_vm_group_bin_1456 = frame (4k)
frame_vm_group_bin_14560 = frame (4k)
frame_vm_group_bin_14561 = frame (4k)
frame_vm_group_bin_14562 = frame (4k)
frame_vm_group_bin_14563 = frame (4k)
frame_vm_group_bin_14564 = frame (4k)
frame_vm_group_bin_14565 = frame (4k)
frame_vm_group_bin_14566 = frame (4k)
frame_vm_group_bin_14567 = frame (4k)
frame_vm_group_bin_14568 = frame (4k)
frame_vm_group_bin_14569 = frame (4k)
frame_vm_group_bin_1457 = frame (4k)
frame_vm_group_bin_14570 = frame (4k)
frame_vm_group_bin_14571 = frame (4k)
frame_vm_group_bin_14572 = frame (4k)
frame_vm_group_bin_14573 = frame (4k)
frame_vm_group_bin_14574 = frame (4k)
frame_vm_group_bin_14575 = frame (4k)
frame_vm_group_bin_14576 = frame (4k)
frame_vm_group_bin_14577 = frame (4k)
frame_vm_group_bin_14578 = frame (4k)
frame_vm_group_bin_14579 = frame (4k)
frame_vm_group_bin_1458 = frame (4k)
frame_vm_group_bin_14580 = frame (4k)
frame_vm_group_bin_14581 = frame (4k)
frame_vm_group_bin_14582 = frame (4k)
frame_vm_group_bin_14583 = frame (4k)
frame_vm_group_bin_14584 = frame (4k)
frame_vm_group_bin_14585 = frame (4k)
frame_vm_group_bin_14586 = frame (4k)
frame_vm_group_bin_14587 = frame (4k)
frame_vm_group_bin_14588 = frame (4k)
frame_vm_group_bin_14589 = frame (4k)
frame_vm_group_bin_1459 = frame (4k)
frame_vm_group_bin_14590 = frame (4k)
frame_vm_group_bin_14591 = frame (4k)
frame_vm_group_bin_14592 = frame (4k)
frame_vm_group_bin_14593 = frame (4k)
frame_vm_group_bin_14594 = frame (4k)
frame_vm_group_bin_14595 = frame (4k)
frame_vm_group_bin_14596 = frame (4k)
frame_vm_group_bin_14597 = frame (4k)
frame_vm_group_bin_14598 = frame (4k)
frame_vm_group_bin_14599 = frame (4k)
frame_vm_group_bin_1460 = frame (4k)
frame_vm_group_bin_14600 = frame (4k)
frame_vm_group_bin_14601 = frame (4k)
frame_vm_group_bin_14602 = frame (4k)
frame_vm_group_bin_14603 = frame (4k)
frame_vm_group_bin_14604 = frame (4k)
frame_vm_group_bin_14605 = frame (4k)
frame_vm_group_bin_14606 = frame (4k)
frame_vm_group_bin_14607 = frame (4k)
frame_vm_group_bin_14608 = frame (4k)
frame_vm_group_bin_14609 = frame (4k)
frame_vm_group_bin_1461 = frame (4k)
frame_vm_group_bin_14610 = frame (4k)
frame_vm_group_bin_14611 = frame (4k)
frame_vm_group_bin_14612 = frame (4k)
frame_vm_group_bin_14613 = frame (4k)
frame_vm_group_bin_14614 = frame (4k)
frame_vm_group_bin_14615 = frame (4k)
frame_vm_group_bin_14616 = frame (4k)
frame_vm_group_bin_14617 = frame (4k)
frame_vm_group_bin_14618 = frame (4k)
frame_vm_group_bin_14619 = frame (4k)
frame_vm_group_bin_1462 = frame (4k)
frame_vm_group_bin_14620 = frame (4k)
frame_vm_group_bin_14621 = frame (4k)
frame_vm_group_bin_14622 = frame (4k)
frame_vm_group_bin_14623 = frame (4k)
frame_vm_group_bin_14624 = frame (4k)
frame_vm_group_bin_14625 = frame (4k)
frame_vm_group_bin_14626 = frame (4k)
frame_vm_group_bin_14627 = frame (4k)
frame_vm_group_bin_14628 = frame (4k)
frame_vm_group_bin_14629 = frame (4k)
frame_vm_group_bin_1463 = frame (4k)
frame_vm_group_bin_14630 = frame (4k)
frame_vm_group_bin_14631 = frame (4k)
frame_vm_group_bin_14632 = frame (4k)
frame_vm_group_bin_14633 = frame (4k)
frame_vm_group_bin_14634 = frame (4k)
frame_vm_group_bin_14635 = frame (4k)
frame_vm_group_bin_14636 = frame (4k)
frame_vm_group_bin_14637 = frame (4k)
frame_vm_group_bin_14638 = frame (4k)
frame_vm_group_bin_14639 = frame (4k)
frame_vm_group_bin_1464 = frame (4k)
frame_vm_group_bin_14640 = frame (4k)
frame_vm_group_bin_14641 = frame (4k)
frame_vm_group_bin_14642 = frame (4k)
frame_vm_group_bin_14643 = frame (4k)
frame_vm_group_bin_14644 = frame (4k)
frame_vm_group_bin_14645 = frame (4k)
frame_vm_group_bin_14646 = frame (4k)
frame_vm_group_bin_14647 = frame (4k)
frame_vm_group_bin_14648 = frame (4k)
frame_vm_group_bin_14649 = frame (4k)
frame_vm_group_bin_1465 = frame (4k)
frame_vm_group_bin_14650 = frame (4k)
frame_vm_group_bin_14651 = frame (4k)
frame_vm_group_bin_14652 = frame (4k)
frame_vm_group_bin_14653 = frame (4k)
frame_vm_group_bin_14654 = frame (4k)
frame_vm_group_bin_14655 = frame (4k)
frame_vm_group_bin_14656 = frame (4k)
frame_vm_group_bin_14657 = frame (4k)
frame_vm_group_bin_14658 = frame (4k)
frame_vm_group_bin_14659 = frame (4k)
frame_vm_group_bin_1466 = frame (4k)
frame_vm_group_bin_14660 = frame (4k)
frame_vm_group_bin_14661 = frame (4k)
frame_vm_group_bin_14662 = frame (4k)
frame_vm_group_bin_14663 = frame (4k)
frame_vm_group_bin_14664 = frame (4k)
frame_vm_group_bin_14665 = frame (4k)
frame_vm_group_bin_14666 = frame (4k)
frame_vm_group_bin_14667 = frame (4k)
frame_vm_group_bin_14668 = frame (4k)
frame_vm_group_bin_14669 = frame (4k)
frame_vm_group_bin_1467 = frame (4k)
frame_vm_group_bin_14670 = frame (4k)
frame_vm_group_bin_14671 = frame (4k)
frame_vm_group_bin_14672 = frame (4k)
frame_vm_group_bin_14673 = frame (4k)
frame_vm_group_bin_14674 = frame (4k)
frame_vm_group_bin_14675 = frame (4k)
frame_vm_group_bin_14676 = frame (4k)
frame_vm_group_bin_14677 = frame (4k)
frame_vm_group_bin_14678 = frame (4k)
frame_vm_group_bin_14679 = frame (4k)
frame_vm_group_bin_1468 = frame (4k)
frame_vm_group_bin_14680 = frame (4k)
frame_vm_group_bin_14681 = frame (4k)
frame_vm_group_bin_14682 = frame (4k)
frame_vm_group_bin_14683 = frame (4k)
frame_vm_group_bin_14684 = frame (4k)
frame_vm_group_bin_14685 = frame (4k)
frame_vm_group_bin_14686 = frame (4k)
frame_vm_group_bin_14687 = frame (4k)
frame_vm_group_bin_14688 = frame (4k)
frame_vm_group_bin_14689 = frame (4k)
frame_vm_group_bin_1469 = frame (4k)
frame_vm_group_bin_14690 = frame (4k)
frame_vm_group_bin_14691 = frame (4k)
frame_vm_group_bin_14692 = frame (4k)
frame_vm_group_bin_14693 = frame (4k)
frame_vm_group_bin_14694 = frame (4k)
frame_vm_group_bin_14695 = frame (4k)
frame_vm_group_bin_14696 = frame (4k)
frame_vm_group_bin_14697 = frame (4k)
frame_vm_group_bin_14698 = frame (4k)
frame_vm_group_bin_14699 = frame (4k)
frame_vm_group_bin_1470 = frame (4k)
frame_vm_group_bin_14700 = frame (4k)
frame_vm_group_bin_14701 = frame (4k)
frame_vm_group_bin_14702 = frame (4k)
frame_vm_group_bin_14703 = frame (4k)
frame_vm_group_bin_14704 = frame (4k)
frame_vm_group_bin_14705 = frame (4k)
frame_vm_group_bin_14706 = frame (4k)
frame_vm_group_bin_14707 = frame (4k)
frame_vm_group_bin_14708 = frame (4k)
frame_vm_group_bin_14709 = frame (4k)
frame_vm_group_bin_1471 = frame (4k)
frame_vm_group_bin_14710 = frame (4k)
frame_vm_group_bin_14711 = frame (4k)
frame_vm_group_bin_14712 = frame (4k)
frame_vm_group_bin_14713 = frame (4k)
frame_vm_group_bin_14714 = frame (4k)
frame_vm_group_bin_14715 = frame (4k)
frame_vm_group_bin_14716 = frame (4k)
frame_vm_group_bin_14717 = frame (4k)
frame_vm_group_bin_14718 = frame (4k)
frame_vm_group_bin_14719 = frame (4k)
frame_vm_group_bin_1472 = frame (4k)
frame_vm_group_bin_14720 = frame (4k)
frame_vm_group_bin_14721 = frame (4k)
frame_vm_group_bin_14722 = frame (4k)
frame_vm_group_bin_14723 = frame (4k)
frame_vm_group_bin_14724 = frame (4k)
frame_vm_group_bin_14725 = frame (4k)
frame_vm_group_bin_14726 = frame (4k)
frame_vm_group_bin_14727 = frame (4k)
frame_vm_group_bin_14728 = frame (4k)
frame_vm_group_bin_14729 = frame (4k)
frame_vm_group_bin_1473 = frame (4k)
frame_vm_group_bin_14730 = frame (4k)
frame_vm_group_bin_14731 = frame (4k)
frame_vm_group_bin_14732 = frame (4k)
frame_vm_group_bin_14733 = frame (4k)
frame_vm_group_bin_14734 = frame (4k)
frame_vm_group_bin_14735 = frame (4k)
frame_vm_group_bin_14736 = frame (4k)
frame_vm_group_bin_14737 = frame (4k)
frame_vm_group_bin_14738 = frame (4k)
frame_vm_group_bin_14739 = frame (4k)
frame_vm_group_bin_1474 = frame (4k)
frame_vm_group_bin_14740 = frame (4k)
frame_vm_group_bin_14741 = frame (4k)
frame_vm_group_bin_14742 = frame (4k)
frame_vm_group_bin_14743 = frame (4k)
frame_vm_group_bin_14744 = frame (4k)
frame_vm_group_bin_14745 = frame (4k)
frame_vm_group_bin_14746 = frame (4k)
frame_vm_group_bin_14747 = frame (4k)
frame_vm_group_bin_14748 = frame (4k)
frame_vm_group_bin_14749 = frame (4k)
frame_vm_group_bin_1475 = frame (4k)
frame_vm_group_bin_14750 = frame (4k)
frame_vm_group_bin_14751 = frame (4k)
frame_vm_group_bin_14752 = frame (4k)
frame_vm_group_bin_14753 = frame (4k)
frame_vm_group_bin_14754 = frame (4k)
frame_vm_group_bin_14755 = frame (4k)
frame_vm_group_bin_14756 = frame (4k)
frame_vm_group_bin_14757 = frame (4k)
frame_vm_group_bin_14758 = frame (4k)
frame_vm_group_bin_14759 = frame (4k)
frame_vm_group_bin_1476 = frame (4k)
frame_vm_group_bin_14760 = frame (4k)
frame_vm_group_bin_14761 = frame (4k)
frame_vm_group_bin_14762 = frame (4k)
frame_vm_group_bin_14763 = frame (4k)
frame_vm_group_bin_14764 = frame (4k)
frame_vm_group_bin_14765 = frame (4k)
frame_vm_group_bin_14766 = frame (4k)
frame_vm_group_bin_14767 = frame (4k)
frame_vm_group_bin_14768 = frame (4k)
frame_vm_group_bin_14769 = frame (4k)
frame_vm_group_bin_1477 = frame (4k)
frame_vm_group_bin_14770 = frame (4k)
frame_vm_group_bin_14771 = frame (4k)
frame_vm_group_bin_14772 = frame (4k)
frame_vm_group_bin_14773 = frame (4k)
frame_vm_group_bin_14774 = frame (4k)
frame_vm_group_bin_14775 = frame (4k)
frame_vm_group_bin_14776 = frame (4k)
frame_vm_group_bin_14777 = frame (4k)
frame_vm_group_bin_14778 = frame (4k)
frame_vm_group_bin_14779 = frame (4k)
frame_vm_group_bin_1478 = frame (4k)
frame_vm_group_bin_14780 = frame (4k)
frame_vm_group_bin_14781 = frame (4k)
frame_vm_group_bin_14782 = frame (4k)
frame_vm_group_bin_14783 = frame (4k)
frame_vm_group_bin_14784 = frame (4k)
frame_vm_group_bin_14785 = frame (4k)
frame_vm_group_bin_14786 = frame (4k)
frame_vm_group_bin_14787 = frame (4k)
frame_vm_group_bin_14788 = frame (4k)
frame_vm_group_bin_14789 = frame (4k)
frame_vm_group_bin_1479 = frame (4k)
frame_vm_group_bin_14790 = frame (4k)
frame_vm_group_bin_14791 = frame (4k)
frame_vm_group_bin_14792 = frame (4k)
frame_vm_group_bin_14793 = frame (4k)
frame_vm_group_bin_14794 = frame (4k)
frame_vm_group_bin_14795 = frame (4k)
frame_vm_group_bin_14796 = frame (4k)
frame_vm_group_bin_14797 = frame (4k)
frame_vm_group_bin_14798 = frame (4k)
frame_vm_group_bin_14799 = frame (4k)
frame_vm_group_bin_1480 = frame (4k)
frame_vm_group_bin_14800 = frame (4k)
frame_vm_group_bin_14801 = frame (4k)
frame_vm_group_bin_14802 = frame (4k)
frame_vm_group_bin_14803 = frame (4k)
frame_vm_group_bin_14804 = frame (4k)
frame_vm_group_bin_14805 = frame (4k)
frame_vm_group_bin_14806 = frame (4k)
frame_vm_group_bin_14807 = frame (4k)
frame_vm_group_bin_14808 = frame (4k)
frame_vm_group_bin_14809 = frame (4k)
frame_vm_group_bin_1481 = frame (4k)
frame_vm_group_bin_14810 = frame (4k)
frame_vm_group_bin_14811 = frame (4k)
frame_vm_group_bin_14812 = frame (4k)
frame_vm_group_bin_14813 = frame (4k)
frame_vm_group_bin_14814 = frame (4k)
frame_vm_group_bin_14815 = frame (4k)
frame_vm_group_bin_14816 = frame (4k)
frame_vm_group_bin_14817 = frame (4k)
frame_vm_group_bin_14818 = frame (4k)
frame_vm_group_bin_14819 = frame (4k)
frame_vm_group_bin_1482 = frame (4k)
frame_vm_group_bin_14820 = frame (4k)
frame_vm_group_bin_14821 = frame (4k)
frame_vm_group_bin_14822 = frame (4k)
frame_vm_group_bin_14823 = frame (4k)
frame_vm_group_bin_14824 = frame (4k)
frame_vm_group_bin_14825 = frame (4k)
frame_vm_group_bin_14826 = frame (4k)
frame_vm_group_bin_14827 = frame (4k)
frame_vm_group_bin_14828 = frame (4k)
frame_vm_group_bin_14829 = frame (4k)
frame_vm_group_bin_1483 = frame (4k)
frame_vm_group_bin_14830 = frame (4k)
frame_vm_group_bin_14831 = frame (4k)
frame_vm_group_bin_14832 = frame (4k)
frame_vm_group_bin_14833 = frame (4k)
frame_vm_group_bin_14834 = frame (4k)
frame_vm_group_bin_14835 = frame (4k)
frame_vm_group_bin_14836 = frame (4k)
frame_vm_group_bin_14837 = frame (4k)
frame_vm_group_bin_14838 = frame (4k)
frame_vm_group_bin_14839 = frame (4k)
frame_vm_group_bin_1484 = frame (4k)
frame_vm_group_bin_14840 = frame (4k)
frame_vm_group_bin_14841 = frame (4k)
frame_vm_group_bin_14842 = frame (4k)
frame_vm_group_bin_14843 = frame (4k)
frame_vm_group_bin_14844 = frame (4k)
frame_vm_group_bin_14845 = frame (4k)
frame_vm_group_bin_14846 = frame (4k)
frame_vm_group_bin_14847 = frame (4k)
frame_vm_group_bin_14848 = frame (4k)
frame_vm_group_bin_14849 = frame (4k)
frame_vm_group_bin_1485 = frame (4k)
frame_vm_group_bin_14850 = frame (4k)
frame_vm_group_bin_14851 = frame (4k)
frame_vm_group_bin_14852 = frame (4k)
frame_vm_group_bin_14853 = frame (4k)
frame_vm_group_bin_14854 = frame (4k)
frame_vm_group_bin_14855 = frame (4k)
frame_vm_group_bin_14856 = frame (4k)
frame_vm_group_bin_14857 = frame (4k)
frame_vm_group_bin_14858 = frame (4k)
frame_vm_group_bin_14859 = frame (4k)
frame_vm_group_bin_1486 = frame (4k)
frame_vm_group_bin_14860 = frame (4k)
frame_vm_group_bin_14861 = frame (4k)
frame_vm_group_bin_14862 = frame (4k)
frame_vm_group_bin_14863 = frame (4k)
frame_vm_group_bin_14864 = frame (4k)
frame_vm_group_bin_14865 = frame (4k)
frame_vm_group_bin_14866 = frame (4k)
frame_vm_group_bin_14867 = frame (4k)
frame_vm_group_bin_14868 = frame (4k)
frame_vm_group_bin_14869 = frame (4k)
frame_vm_group_bin_1487 = frame (4k)
frame_vm_group_bin_14870 = frame (4k)
frame_vm_group_bin_14871 = frame (4k)
frame_vm_group_bin_14872 = frame (4k)
frame_vm_group_bin_14873 = frame (4k)
frame_vm_group_bin_14874 = frame (4k)
frame_vm_group_bin_14875 = frame (4k)
frame_vm_group_bin_14876 = frame (4k)
frame_vm_group_bin_14877 = frame (4k)
frame_vm_group_bin_14878 = frame (4k)
frame_vm_group_bin_14879 = frame (4k)
frame_vm_group_bin_1488 = frame (4k)
frame_vm_group_bin_14880 = frame (4k)
frame_vm_group_bin_14881 = frame (4k)
frame_vm_group_bin_14882 = frame (4k)
frame_vm_group_bin_14883 = frame (4k)
frame_vm_group_bin_14884 = frame (4k)
frame_vm_group_bin_14885 = frame (4k)
frame_vm_group_bin_14886 = frame (4k)
frame_vm_group_bin_14887 = frame (4k)
frame_vm_group_bin_14888 = frame (4k)
frame_vm_group_bin_14889 = frame (4k)
frame_vm_group_bin_1489 = frame (4k)
frame_vm_group_bin_14890 = frame (4k)
frame_vm_group_bin_14891 = frame (4k)
frame_vm_group_bin_14892 = frame (4k)
frame_vm_group_bin_14893 = frame (4k)
frame_vm_group_bin_14894 = frame (4k)
frame_vm_group_bin_14895 = frame (4k)
frame_vm_group_bin_14896 = frame (4k)
frame_vm_group_bin_14897 = frame (4k)
frame_vm_group_bin_14898 = frame (4k)
frame_vm_group_bin_14899 = frame (4k)
frame_vm_group_bin_1490 = frame (4k)
frame_vm_group_bin_14900 = frame (4k)
frame_vm_group_bin_14901 = frame (4k)
frame_vm_group_bin_14902 = frame (4k)
frame_vm_group_bin_14903 = frame (4k)
frame_vm_group_bin_14904 = frame (4k)
frame_vm_group_bin_14905 = frame (4k)
frame_vm_group_bin_14906 = frame (4k)
frame_vm_group_bin_14907 = frame (4k)
frame_vm_group_bin_14908 = frame (4k)
frame_vm_group_bin_14909 = frame (4k)
frame_vm_group_bin_1491 = frame (4k)
frame_vm_group_bin_14910 = frame (4k)
frame_vm_group_bin_14911 = frame (4k)
frame_vm_group_bin_14912 = frame (4k)
frame_vm_group_bin_14913 = frame (4k)
frame_vm_group_bin_14914 = frame (4k)
frame_vm_group_bin_14915 = frame (4k)
frame_vm_group_bin_14916 = frame (4k)
frame_vm_group_bin_14917 = frame (4k)
frame_vm_group_bin_14918 = frame (4k)
frame_vm_group_bin_14919 = frame (4k)
frame_vm_group_bin_1492 = frame (4k)
frame_vm_group_bin_14920 = frame (4k)
frame_vm_group_bin_14921 = frame (4k)
frame_vm_group_bin_14922 = frame (4k)
frame_vm_group_bin_14923 = frame (4k)
frame_vm_group_bin_14924 = frame (4k)
frame_vm_group_bin_14925 = frame (4k)
frame_vm_group_bin_14926 = frame (4k)
frame_vm_group_bin_14927 = frame (4k)
frame_vm_group_bin_14928 = frame (4k)
frame_vm_group_bin_14929 = frame (4k)
frame_vm_group_bin_1493 = frame (4k)
frame_vm_group_bin_14930 = frame (4k)
frame_vm_group_bin_14931 = frame (4k)
frame_vm_group_bin_14932 = frame (4k)
frame_vm_group_bin_14933 = frame (4k)
frame_vm_group_bin_14934 = frame (4k)
frame_vm_group_bin_14935 = frame (4k)
frame_vm_group_bin_14936 = frame (4k)
frame_vm_group_bin_14937 = frame (4k)
frame_vm_group_bin_14938 = frame (4k)
frame_vm_group_bin_14939 = frame (4k)
frame_vm_group_bin_1494 = frame (4k)
frame_vm_group_bin_14940 = frame (4k)
frame_vm_group_bin_14941 = frame (4k)
frame_vm_group_bin_14942 = frame (4k)
frame_vm_group_bin_14943 = frame (4k)
frame_vm_group_bin_14944 = frame (4k)
frame_vm_group_bin_14945 = frame (4k)
frame_vm_group_bin_14946 = frame (4k)
frame_vm_group_bin_14947 = frame (4k)
frame_vm_group_bin_14948 = frame (4k)
frame_vm_group_bin_14949 = frame (4k)
frame_vm_group_bin_1495 = frame (4k)
frame_vm_group_bin_14950 = frame (4k)
frame_vm_group_bin_14951 = frame (4k)
frame_vm_group_bin_14952 = frame (4k)
frame_vm_group_bin_14953 = frame (4k)
frame_vm_group_bin_14954 = frame (4k)
frame_vm_group_bin_14955 = frame (4k)
frame_vm_group_bin_14956 = frame (4k)
frame_vm_group_bin_14957 = frame (4k)
frame_vm_group_bin_14958 = frame (4k)
frame_vm_group_bin_14959 = frame (4k)
frame_vm_group_bin_1496 = frame (4k)
frame_vm_group_bin_14960 = frame (4k)
frame_vm_group_bin_14961 = frame (4k)
frame_vm_group_bin_14962 = frame (4k)
frame_vm_group_bin_14963 = frame (4k)
frame_vm_group_bin_14964 = frame (4k)
frame_vm_group_bin_14965 = frame (4k)
frame_vm_group_bin_14966 = frame (4k)
frame_vm_group_bin_14967 = frame (4k)
frame_vm_group_bin_14968 = frame (4k)
frame_vm_group_bin_14969 = frame (4k)
frame_vm_group_bin_1497 = frame (4k)
frame_vm_group_bin_14970 = frame (4k)
frame_vm_group_bin_14971 = frame (4k)
frame_vm_group_bin_14972 = frame (4k)
frame_vm_group_bin_14973 = frame (4k)
frame_vm_group_bin_14974 = frame (4k)
frame_vm_group_bin_14975 = frame (4k)
frame_vm_group_bin_14976 = frame (4k)
frame_vm_group_bin_14977 = frame (4k)
frame_vm_group_bin_14978 = frame (4k)
frame_vm_group_bin_14979 = frame (4k)
frame_vm_group_bin_1498 = frame (4k)
frame_vm_group_bin_14980 = frame (4k)
frame_vm_group_bin_14981 = frame (4k)
frame_vm_group_bin_14982 = frame (4k)
frame_vm_group_bin_14983 = frame (4k)
frame_vm_group_bin_14984 = frame (4k)
frame_vm_group_bin_14985 = frame (4k)
frame_vm_group_bin_14986 = frame (4k)
frame_vm_group_bin_14987 = frame (4k)
frame_vm_group_bin_14988 = frame (4k)
frame_vm_group_bin_14989 = frame (4k)
frame_vm_group_bin_1499 = frame (4k)
frame_vm_group_bin_14990 = frame (4k)
frame_vm_group_bin_14991 = frame (4k)
frame_vm_group_bin_14992 = frame (4k)
frame_vm_group_bin_14993 = frame (4k)
frame_vm_group_bin_14994 = frame (4k)
frame_vm_group_bin_14995 = frame (4k)
frame_vm_group_bin_14996 = frame (4k)
frame_vm_group_bin_14997 = frame (4k)
frame_vm_group_bin_14998 = frame (4k)
frame_vm_group_bin_14999 = frame (4k)
frame_vm_group_bin_1500 = frame (4k)
frame_vm_group_bin_15000 = frame (4k)
frame_vm_group_bin_15001 = frame (4k)
frame_vm_group_bin_15002 = frame (4k)
frame_vm_group_bin_15003 = frame (4k)
frame_vm_group_bin_15004 = frame (4k)
frame_vm_group_bin_15005 = frame (4k)
frame_vm_group_bin_15006 = frame (4k)
frame_vm_group_bin_15007 = frame (4k)
frame_vm_group_bin_15008 = frame (4k)
frame_vm_group_bin_15009 = frame (4k)
frame_vm_group_bin_1501 = frame (4k)
frame_vm_group_bin_15010 = frame (4k)
frame_vm_group_bin_15011 = frame (4k)
frame_vm_group_bin_15012 = frame (4k)
frame_vm_group_bin_15013 = frame (4k)
frame_vm_group_bin_15014 = frame (4k)
frame_vm_group_bin_15015 = frame (4k)
frame_vm_group_bin_15016 = frame (4k)
frame_vm_group_bin_15017 = frame (4k)
frame_vm_group_bin_15018 = frame (4k)
frame_vm_group_bin_15019 = frame (4k)
frame_vm_group_bin_1502 = frame (4k)
frame_vm_group_bin_15020 = frame (4k)
frame_vm_group_bin_15021 = frame (4k)
frame_vm_group_bin_15022 = frame (4k)
frame_vm_group_bin_15023 = frame (4k)
frame_vm_group_bin_15024 = frame (4k)
frame_vm_group_bin_15025 = frame (4k)
frame_vm_group_bin_15026 = frame (4k)
frame_vm_group_bin_15027 = frame (4k)
frame_vm_group_bin_15028 = frame (4k)
frame_vm_group_bin_15029 = frame (4k)
frame_vm_group_bin_1503 = frame (4k)
frame_vm_group_bin_15030 = frame (4k)
frame_vm_group_bin_15031 = frame (4k)
frame_vm_group_bin_15032 = frame (4k)
frame_vm_group_bin_15033 = frame (4k)
frame_vm_group_bin_15034 = frame (4k)
frame_vm_group_bin_15035 = frame (4k)
frame_vm_group_bin_15036 = frame (4k)
frame_vm_group_bin_15037 = frame (4k)
frame_vm_group_bin_15038 = frame (4k)
frame_vm_group_bin_15039 = frame (4k)
frame_vm_group_bin_1504 = frame (4k)
frame_vm_group_bin_15040 = frame (4k)
frame_vm_group_bin_15041 = frame (4k)
frame_vm_group_bin_15042 = frame (4k)
frame_vm_group_bin_15043 = frame (4k)
frame_vm_group_bin_15044 = frame (4k)
frame_vm_group_bin_15045 = frame (4k)
frame_vm_group_bin_15046 = frame (4k)
frame_vm_group_bin_15047 = frame (4k)
frame_vm_group_bin_15048 = frame (4k)
frame_vm_group_bin_15049 = frame (4k)
frame_vm_group_bin_1505 = frame (4k)
frame_vm_group_bin_15050 = frame (4k)
frame_vm_group_bin_15051 = frame (4k)
frame_vm_group_bin_15052 = frame (4k)
frame_vm_group_bin_15053 = frame (4k)
frame_vm_group_bin_15054 = frame (4k)
frame_vm_group_bin_15055 = frame (4k)
frame_vm_group_bin_15056 = frame (4k)
frame_vm_group_bin_15057 = frame (4k)
frame_vm_group_bin_15058 = frame (4k)
frame_vm_group_bin_15059 = frame (4k)
frame_vm_group_bin_1506 = frame (4k)
frame_vm_group_bin_15060 = frame (4k)
frame_vm_group_bin_15061 = frame (4k)
frame_vm_group_bin_15062 = frame (4k)
frame_vm_group_bin_15063 = frame (4k)
frame_vm_group_bin_15064 = frame (4k)
frame_vm_group_bin_15065 = frame (4k)
frame_vm_group_bin_15066 = frame (4k)
frame_vm_group_bin_15067 = frame (4k)
frame_vm_group_bin_15068 = frame (4k)
frame_vm_group_bin_15069 = frame (4k)
frame_vm_group_bin_1507 = frame (4k)
frame_vm_group_bin_15070 = frame (4k)
frame_vm_group_bin_15071 = frame (4k)
frame_vm_group_bin_15072 = frame (4k)
frame_vm_group_bin_15073 = frame (4k)
frame_vm_group_bin_15074 = frame (4k)
frame_vm_group_bin_15075 = frame (4k)
frame_vm_group_bin_15076 = frame (4k)
frame_vm_group_bin_15077 = frame (4k)
frame_vm_group_bin_15078 = frame (4k)
frame_vm_group_bin_15079 = frame (4k)
frame_vm_group_bin_1508 = frame (4k)
frame_vm_group_bin_15080 = frame (4k)
frame_vm_group_bin_15081 = frame (4k)
frame_vm_group_bin_15082 = frame (4k)
frame_vm_group_bin_15083 = frame (4k)
frame_vm_group_bin_15084 = frame (4k)
frame_vm_group_bin_15085 = frame (4k)
frame_vm_group_bin_15086 = frame (4k)
frame_vm_group_bin_15087 = frame (4k)
frame_vm_group_bin_15088 = frame (4k)
frame_vm_group_bin_15089 = frame (4k)
frame_vm_group_bin_1509 = frame (4k)
frame_vm_group_bin_15090 = frame (4k)
frame_vm_group_bin_15091 = frame (4k)
frame_vm_group_bin_15092 = frame (4k)
frame_vm_group_bin_15093 = frame (4k)
frame_vm_group_bin_15094 = frame (4k)
frame_vm_group_bin_15095 = frame (4k)
frame_vm_group_bin_15096 = frame (4k)
frame_vm_group_bin_15097 = frame (4k)
frame_vm_group_bin_15098 = frame (4k)
frame_vm_group_bin_15099 = frame (4k)
frame_vm_group_bin_1510 = frame (4k)
frame_vm_group_bin_15100 = frame (4k)
frame_vm_group_bin_15101 = frame (4k)
frame_vm_group_bin_15102 = frame (4k)
frame_vm_group_bin_15103 = frame (4k)
frame_vm_group_bin_15104 = frame (4k)
frame_vm_group_bin_15105 = frame (4k)
frame_vm_group_bin_15106 = frame (4k)
frame_vm_group_bin_15107 = frame (4k)
frame_vm_group_bin_15108 = frame (4k)
frame_vm_group_bin_15109 = frame (4k)
frame_vm_group_bin_1511 = frame (4k)
frame_vm_group_bin_15110 = frame (4k)
frame_vm_group_bin_15111 = frame (4k)
frame_vm_group_bin_15112 = frame (4k)
frame_vm_group_bin_15113 = frame (4k)
frame_vm_group_bin_15114 = frame (4k)
frame_vm_group_bin_15115 = frame (4k)
frame_vm_group_bin_15116 = frame (4k)
frame_vm_group_bin_15117 = frame (4k)
frame_vm_group_bin_15118 = frame (4k)
frame_vm_group_bin_15119 = frame (4k)
frame_vm_group_bin_1512 = frame (4k)
frame_vm_group_bin_15120 = frame (4k)
frame_vm_group_bin_15121 = frame (4k)
frame_vm_group_bin_15122 = frame (4k)
frame_vm_group_bin_15123 = frame (4k)
frame_vm_group_bin_15124 = frame (4k)
frame_vm_group_bin_15125 = frame (4k)
frame_vm_group_bin_15126 = frame (4k)
frame_vm_group_bin_15127 = frame (4k)
frame_vm_group_bin_15128 = frame (4k)
frame_vm_group_bin_15129 = frame (4k)
frame_vm_group_bin_1513 = frame (4k)
frame_vm_group_bin_15130 = frame (4k)
frame_vm_group_bin_15131 = frame (4k)
frame_vm_group_bin_15132 = frame (4k)
frame_vm_group_bin_15133 = frame (4k)
frame_vm_group_bin_15134 = frame (4k)
frame_vm_group_bin_15135 = frame (4k)
frame_vm_group_bin_15136 = frame (4k)
frame_vm_group_bin_15137 = frame (4k)
frame_vm_group_bin_15138 = frame (4k)
frame_vm_group_bin_15139 = frame (4k)
frame_vm_group_bin_1514 = frame (4k)
frame_vm_group_bin_15140 = frame (4k)
frame_vm_group_bin_15141 = frame (4k)
frame_vm_group_bin_15142 = frame (4k)
frame_vm_group_bin_15143 = frame (4k)
frame_vm_group_bin_15144 = frame (4k)
frame_vm_group_bin_15145 = frame (4k)
frame_vm_group_bin_15146 = frame (4k)
frame_vm_group_bin_15147 = frame (4k)
frame_vm_group_bin_15148 = frame (4k)
frame_vm_group_bin_15149 = frame (4k)
frame_vm_group_bin_1515 = frame (4k)
frame_vm_group_bin_15150 = frame (4k)
frame_vm_group_bin_15151 = frame (4k)
frame_vm_group_bin_15152 = frame (4k)
frame_vm_group_bin_15153 = frame (4k)
frame_vm_group_bin_15154 = frame (4k)
frame_vm_group_bin_15155 = frame (4k)
frame_vm_group_bin_15156 = frame (4k)
frame_vm_group_bin_15157 = frame (4k)
frame_vm_group_bin_15158 = frame (4k)
frame_vm_group_bin_15159 = frame (4k)
frame_vm_group_bin_1516 = frame (4k)
frame_vm_group_bin_15160 = frame (4k)
frame_vm_group_bin_15161 = frame (4k)
frame_vm_group_bin_15162 = frame (4k)
frame_vm_group_bin_15163 = frame (4k)
frame_vm_group_bin_15164 = frame (4k)
frame_vm_group_bin_15165 = frame (4k)
frame_vm_group_bin_15166 = frame (4k)
frame_vm_group_bin_15167 = frame (4k)
frame_vm_group_bin_15168 = frame (4k)
frame_vm_group_bin_15169 = frame (4k)
frame_vm_group_bin_1517 = frame (4k)
frame_vm_group_bin_15170 = frame (4k)
frame_vm_group_bin_15171 = frame (4k)
frame_vm_group_bin_15172 = frame (4k)
frame_vm_group_bin_15173 = frame (4k)
frame_vm_group_bin_15174 = frame (4k)
frame_vm_group_bin_15175 = frame (4k)
frame_vm_group_bin_15176 = frame (4k)
frame_vm_group_bin_15177 = frame (4k)
frame_vm_group_bin_15178 = frame (4k)
frame_vm_group_bin_15179 = frame (4k)
frame_vm_group_bin_1518 = frame (4k)
frame_vm_group_bin_15180 = frame (4k)
frame_vm_group_bin_15181 = frame (4k)
frame_vm_group_bin_15182 = frame (4k)
frame_vm_group_bin_15183 = frame (4k)
frame_vm_group_bin_15184 = frame (4k)
frame_vm_group_bin_15185 = frame (4k)
frame_vm_group_bin_15186 = frame (4k)
frame_vm_group_bin_15187 = frame (4k)
frame_vm_group_bin_15188 = frame (4k)
frame_vm_group_bin_15189 = frame (4k)
frame_vm_group_bin_1519 = frame (4k)
frame_vm_group_bin_15190 = frame (4k)
frame_vm_group_bin_15191 = frame (4k)
frame_vm_group_bin_15192 = frame (4k)
frame_vm_group_bin_15193 = frame (4k)
frame_vm_group_bin_15194 = frame (4k)
frame_vm_group_bin_15195 = frame (4k)
frame_vm_group_bin_15196 = frame (4k)
frame_vm_group_bin_15197 = frame (4k)
frame_vm_group_bin_15198 = frame (4k)
frame_vm_group_bin_15199 = frame (4k)
frame_vm_group_bin_1520 = frame (4k)
frame_vm_group_bin_15200 = frame (4k)
frame_vm_group_bin_15201 = frame (4k)
frame_vm_group_bin_15202 = frame (4k)
frame_vm_group_bin_15203 = frame (4k)
frame_vm_group_bin_15204 = frame (4k)
frame_vm_group_bin_15205 = frame (4k)
frame_vm_group_bin_15206 = frame (4k)
frame_vm_group_bin_15207 = frame (4k)
frame_vm_group_bin_15208 = frame (4k)
frame_vm_group_bin_15209 = frame (4k)
frame_vm_group_bin_1521 = frame (4k)
frame_vm_group_bin_15210 = frame (4k)
frame_vm_group_bin_15211 = frame (4k)
frame_vm_group_bin_15212 = frame (4k)
frame_vm_group_bin_15213 = frame (4k)
frame_vm_group_bin_15214 = frame (4k)
frame_vm_group_bin_15215 = frame (4k)
frame_vm_group_bin_15216 = frame (4k)
frame_vm_group_bin_15217 = frame (4k)
frame_vm_group_bin_15218 = frame (4k)
frame_vm_group_bin_15219 = frame (4k)
frame_vm_group_bin_1522 = frame (4k)
frame_vm_group_bin_15220 = frame (4k)
frame_vm_group_bin_15221 = frame (4k)
frame_vm_group_bin_15222 = frame (4k)
frame_vm_group_bin_15223 = frame (4k)
frame_vm_group_bin_15224 = frame (4k)
frame_vm_group_bin_15225 = frame (4k)
frame_vm_group_bin_15226 = frame (4k)
frame_vm_group_bin_15227 = frame (4k)
frame_vm_group_bin_15228 = frame (4k)
frame_vm_group_bin_15229 = frame (4k)
frame_vm_group_bin_1523 = frame (4k)
frame_vm_group_bin_15230 = frame (4k)
frame_vm_group_bin_15231 = frame (4k)
frame_vm_group_bin_15232 = frame (4k)
frame_vm_group_bin_15233 = frame (4k)
frame_vm_group_bin_15234 = frame (4k)
frame_vm_group_bin_15235 = frame (4k)
frame_vm_group_bin_15236 = frame (4k)
frame_vm_group_bin_15237 = frame (4k)
frame_vm_group_bin_15238 = frame (4k)
frame_vm_group_bin_15239 = frame (4k)
frame_vm_group_bin_1524 = frame (4k)
frame_vm_group_bin_15240 = frame (4k)
frame_vm_group_bin_15241 = frame (4k)
frame_vm_group_bin_15242 = frame (4k)
frame_vm_group_bin_15243 = frame (4k)
frame_vm_group_bin_15244 = frame (4k)
frame_vm_group_bin_15245 = frame (4k)
frame_vm_group_bin_15246 = frame (4k)
frame_vm_group_bin_15247 = frame (4k)
frame_vm_group_bin_15248 = frame (4k)
frame_vm_group_bin_15249 = frame (4k)
frame_vm_group_bin_1525 = frame (4k)
frame_vm_group_bin_15250 = frame (4k)
frame_vm_group_bin_15251 = frame (4k)
frame_vm_group_bin_15252 = frame (4k)
frame_vm_group_bin_15253 = frame (4k)
frame_vm_group_bin_15254 = frame (4k)
frame_vm_group_bin_15255 = frame (4k)
frame_vm_group_bin_15256 = frame (4k)
frame_vm_group_bin_15257 = frame (4k)
frame_vm_group_bin_15258 = frame (4k)
frame_vm_group_bin_15259 = frame (4k)
frame_vm_group_bin_1526 = frame (4k)
frame_vm_group_bin_15260 = frame (4k)
frame_vm_group_bin_15261 = frame (4k)
frame_vm_group_bin_15262 = frame (4k)
frame_vm_group_bin_15263 = frame (4k)
frame_vm_group_bin_15264 = frame (4k)
frame_vm_group_bin_15265 = frame (4k)
frame_vm_group_bin_15266 = frame (4k)
frame_vm_group_bin_15267 = frame (4k)
frame_vm_group_bin_15268 = frame (4k)
frame_vm_group_bin_15269 = frame (4k)
frame_vm_group_bin_1527 = frame (4k)
frame_vm_group_bin_15270 = frame (4k)
frame_vm_group_bin_15271 = frame (4k)
frame_vm_group_bin_15272 = frame (4k)
frame_vm_group_bin_15273 = frame (4k)
frame_vm_group_bin_15274 = frame (4k)
frame_vm_group_bin_15275 = frame (4k)
frame_vm_group_bin_15276 = frame (4k)
frame_vm_group_bin_15277 = frame (4k)
frame_vm_group_bin_15278 = frame (4k)
frame_vm_group_bin_15279 = frame (4k)
frame_vm_group_bin_1528 = frame (4k)
frame_vm_group_bin_15280 = frame (4k)
frame_vm_group_bin_15281 = frame (4k)
frame_vm_group_bin_15282 = frame (4k)
frame_vm_group_bin_15283 = frame (4k)
frame_vm_group_bin_15284 = frame (4k)
frame_vm_group_bin_15285 = frame (4k)
frame_vm_group_bin_15286 = frame (4k)
frame_vm_group_bin_15287 = frame (4k)
frame_vm_group_bin_15288 = frame (4k)
frame_vm_group_bin_15289 = frame (4k)
frame_vm_group_bin_1529 = frame (4k)
frame_vm_group_bin_15290 = frame (4k)
frame_vm_group_bin_15291 = frame (4k)
frame_vm_group_bin_15292 = frame (4k)
frame_vm_group_bin_15293 = frame (4k)
frame_vm_group_bin_15294 = frame (4k)
frame_vm_group_bin_15295 = frame (4k)
frame_vm_group_bin_15296 = frame (4k)
frame_vm_group_bin_15297 = frame (4k)
frame_vm_group_bin_15298 = frame (4k)
frame_vm_group_bin_15299 = frame (4k)
frame_vm_group_bin_1530 = frame (4k)
frame_vm_group_bin_15300 = frame (4k)
frame_vm_group_bin_15301 = frame (4k)
frame_vm_group_bin_15302 = frame (4k)
frame_vm_group_bin_15303 = frame (4k)
frame_vm_group_bin_15304 = frame (4k)
frame_vm_group_bin_15305 = frame (4k)
frame_vm_group_bin_15306 = frame (4k)
frame_vm_group_bin_15307 = frame (4k)
frame_vm_group_bin_15308 = frame (4k)
frame_vm_group_bin_15309 = frame (4k)
frame_vm_group_bin_1531 = frame (4k)
frame_vm_group_bin_15310 = frame (4k)
frame_vm_group_bin_15311 = frame (4k)
frame_vm_group_bin_15312 = frame (4k)
frame_vm_group_bin_15313 = frame (4k)
frame_vm_group_bin_15314 = frame (4k)
frame_vm_group_bin_15315 = frame (4k)
frame_vm_group_bin_15316 = frame (4k)
frame_vm_group_bin_15317 = frame (4k)
frame_vm_group_bin_15318 = frame (4k)
frame_vm_group_bin_15319 = frame (4k)
frame_vm_group_bin_1532 = frame (4k)
frame_vm_group_bin_15320 = frame (4k)
frame_vm_group_bin_15321 = frame (4k)
frame_vm_group_bin_15322 = frame (4k)
frame_vm_group_bin_15323 = frame (4k)
frame_vm_group_bin_15324 = frame (4k)
frame_vm_group_bin_15325 = frame (4k)
frame_vm_group_bin_15326 = frame (4k)
frame_vm_group_bin_15327 = frame (4k)
frame_vm_group_bin_15328 = frame (4k)
frame_vm_group_bin_15329 = frame (4k)
frame_vm_group_bin_1533 = frame (4k)
frame_vm_group_bin_15330 = frame (4k)
frame_vm_group_bin_15331 = frame (4k)
frame_vm_group_bin_15332 = frame (4k)
frame_vm_group_bin_15333 = frame (4k)
frame_vm_group_bin_15334 = frame (4k)
frame_vm_group_bin_15335 = frame (4k)
frame_vm_group_bin_15336 = frame (4k)
frame_vm_group_bin_15337 = frame (4k)
frame_vm_group_bin_15338 = frame (4k)
frame_vm_group_bin_15339 = frame (4k)
frame_vm_group_bin_1534 = frame (4k)
frame_vm_group_bin_15340 = frame (4k)
frame_vm_group_bin_15341 = frame (4k)
frame_vm_group_bin_15342 = frame (4k)
frame_vm_group_bin_15343 = frame (4k)
frame_vm_group_bin_15344 = frame (4k)
frame_vm_group_bin_15345 = frame (4k)
frame_vm_group_bin_15346 = frame (4k)
frame_vm_group_bin_15347 = frame (4k)
frame_vm_group_bin_15348 = frame (4k)
frame_vm_group_bin_15349 = frame (4k)
frame_vm_group_bin_1535 = frame (4k)
frame_vm_group_bin_15350 = frame (4k)
frame_vm_group_bin_15351 = frame (4k)
frame_vm_group_bin_15352 = frame (4k)
frame_vm_group_bin_15353 = frame (4k)
frame_vm_group_bin_15354 = frame (4k)
frame_vm_group_bin_15355 = frame (4k)
frame_vm_group_bin_15356 = frame (4k)
frame_vm_group_bin_15357 = frame (4k)
frame_vm_group_bin_15358 = frame (4k)
frame_vm_group_bin_15359 = frame (4k)
frame_vm_group_bin_1536 = frame (4k)
frame_vm_group_bin_15360 = frame (4k)
frame_vm_group_bin_15361 = frame (4k)
frame_vm_group_bin_15362 = frame (4k)
frame_vm_group_bin_15363 = frame (4k)
frame_vm_group_bin_15364 = frame (4k)
frame_vm_group_bin_15365 = frame (4k)
frame_vm_group_bin_15366 = frame (4k)
frame_vm_group_bin_15367 = frame (4k)
frame_vm_group_bin_15368 = frame (4k)
frame_vm_group_bin_15369 = frame (4k)
frame_vm_group_bin_1537 = frame (4k)
frame_vm_group_bin_15370 = frame (4k)
frame_vm_group_bin_15371 = frame (4k)
frame_vm_group_bin_15372 = frame (4k)
frame_vm_group_bin_15373 = frame (4k)
frame_vm_group_bin_15374 = frame (4k)
frame_vm_group_bin_15375 = frame (4k)
frame_vm_group_bin_15376 = frame (4k)
frame_vm_group_bin_15377 = frame (4k)
frame_vm_group_bin_15378 = frame (4k)
frame_vm_group_bin_15379 = frame (4k)
frame_vm_group_bin_1538 = frame (4k)
frame_vm_group_bin_15380 = frame (4k)
frame_vm_group_bin_15381 = frame (4k)
frame_vm_group_bin_15382 = frame (4k)
frame_vm_group_bin_15383 = frame (4k)
frame_vm_group_bin_15384 = frame (4k)
frame_vm_group_bin_15385 = frame (4k)
frame_vm_group_bin_15386 = frame (4k)
frame_vm_group_bin_15387 = frame (4k)
frame_vm_group_bin_15388 = frame (4k)
frame_vm_group_bin_15389 = frame (4k)
frame_vm_group_bin_1539 = frame (4k)
frame_vm_group_bin_15390 = frame (4k)
frame_vm_group_bin_15391 = frame (4k)
frame_vm_group_bin_15392 = frame (4k)
frame_vm_group_bin_15393 = frame (4k)
frame_vm_group_bin_15394 = frame (4k)
frame_vm_group_bin_15395 = frame (4k)
frame_vm_group_bin_15396 = frame (4k)
frame_vm_group_bin_15397 = frame (4k)
frame_vm_group_bin_15398 = frame (4k)
frame_vm_group_bin_15399 = frame (4k)
frame_vm_group_bin_1540 = frame (4k)
frame_vm_group_bin_15400 = frame (4k)
frame_vm_group_bin_15401 = frame (4k)
frame_vm_group_bin_15402 = frame (4k)
frame_vm_group_bin_15403 = frame (4k)
frame_vm_group_bin_15404 = frame (4k)
frame_vm_group_bin_15405 = frame (4k)
frame_vm_group_bin_15406 = frame (4k)
frame_vm_group_bin_15407 = frame (4k)
frame_vm_group_bin_15408 = frame (4k)
frame_vm_group_bin_15409 = frame (4k)
frame_vm_group_bin_1541 = frame (4k)
frame_vm_group_bin_15410 = frame (4k)
frame_vm_group_bin_15411 = frame (4k)
frame_vm_group_bin_15412 = frame (4k)
frame_vm_group_bin_15413 = frame (4k)
frame_vm_group_bin_15414 = frame (4k)
frame_vm_group_bin_15415 = frame (4k)
frame_vm_group_bin_15416 = frame (4k)
frame_vm_group_bin_15417 = frame (4k)
frame_vm_group_bin_15418 = frame (4k)
frame_vm_group_bin_15419 = frame (4k)
frame_vm_group_bin_1542 = frame (4k)
frame_vm_group_bin_15420 = frame (4k)
frame_vm_group_bin_15421 = frame (4k)
frame_vm_group_bin_15422 = frame (4k)
frame_vm_group_bin_15423 = frame (4k)
frame_vm_group_bin_15424 = frame (4k)
frame_vm_group_bin_15425 = frame (4k)
frame_vm_group_bin_15426 = frame (4k)
frame_vm_group_bin_15427 = frame (4k)
frame_vm_group_bin_15428 = frame (4k)
frame_vm_group_bin_15429 = frame (4k)
frame_vm_group_bin_1543 = frame (4k)
frame_vm_group_bin_15430 = frame (4k)
frame_vm_group_bin_15431 = frame (4k)
frame_vm_group_bin_15432 = frame (4k)
frame_vm_group_bin_15433 = frame (4k)
frame_vm_group_bin_15434 = frame (4k)
frame_vm_group_bin_15435 = frame (4k)
frame_vm_group_bin_15436 = frame (4k)
frame_vm_group_bin_15437 = frame (4k)
frame_vm_group_bin_15438 = frame (4k)
frame_vm_group_bin_15439 = frame (4k)
frame_vm_group_bin_1544 = frame (4k)
frame_vm_group_bin_15440 = frame (4k)
frame_vm_group_bin_15441 = frame (4k)
frame_vm_group_bin_15442 = frame (4k)
frame_vm_group_bin_15443 = frame (4k)
frame_vm_group_bin_15444 = frame (4k)
frame_vm_group_bin_15445 = frame (4k)
frame_vm_group_bin_15446 = frame (4k)
frame_vm_group_bin_15447 = frame (4k)
frame_vm_group_bin_15448 = frame (4k)
frame_vm_group_bin_15449 = frame (4k)
frame_vm_group_bin_1545 = frame (4k)
frame_vm_group_bin_15450 = frame (4k)
frame_vm_group_bin_15451 = frame (4k)
frame_vm_group_bin_15452 = frame (4k)
frame_vm_group_bin_15453 = frame (4k)
frame_vm_group_bin_15454 = frame (4k)
frame_vm_group_bin_15455 = frame (4k)
frame_vm_group_bin_15456 = frame (4k)
frame_vm_group_bin_15457 = frame (4k)
frame_vm_group_bin_15458 = frame (4k)
frame_vm_group_bin_15459 = frame (4k)
frame_vm_group_bin_1546 = frame (4k)
frame_vm_group_bin_15460 = frame (4k)
frame_vm_group_bin_15461 = frame (4k)
frame_vm_group_bin_15462 = frame (4k)
frame_vm_group_bin_15463 = frame (4k)
frame_vm_group_bin_15464 = frame (4k)
frame_vm_group_bin_15465 = frame (4k)
frame_vm_group_bin_15466 = frame (4k)
frame_vm_group_bin_15467 = frame (4k)
frame_vm_group_bin_15468 = frame (4k)
frame_vm_group_bin_15469 = frame (4k)
frame_vm_group_bin_1547 = frame (4k)
frame_vm_group_bin_15470 = frame (4k)
frame_vm_group_bin_15471 = frame (4k)
frame_vm_group_bin_15472 = frame (4k)
frame_vm_group_bin_15473 = frame (4k)
frame_vm_group_bin_15474 = frame (4k)
frame_vm_group_bin_15475 = frame (4k)
frame_vm_group_bin_15476 = frame (4k)
frame_vm_group_bin_15477 = frame (4k)
frame_vm_group_bin_15478 = frame (4k)
frame_vm_group_bin_15479 = frame (4k)
frame_vm_group_bin_1548 = frame (4k)
frame_vm_group_bin_15480 = frame (4k)
frame_vm_group_bin_15481 = frame (4k)
frame_vm_group_bin_15482 = frame (4k)
frame_vm_group_bin_15483 = frame (4k)
frame_vm_group_bin_15484 = frame (4k)
frame_vm_group_bin_15485 = frame (4k)
frame_vm_group_bin_15486 = frame (4k)
frame_vm_group_bin_15487 = frame (4k)
frame_vm_group_bin_15488 = frame (4k)
frame_vm_group_bin_15489 = frame (4k)
frame_vm_group_bin_1549 = frame (4k)
frame_vm_group_bin_15490 = frame (4k)
frame_vm_group_bin_15491 = frame (4k)
frame_vm_group_bin_15492 = frame (4k)
frame_vm_group_bin_15493 = frame (4k)
frame_vm_group_bin_15494 = frame (4k)
frame_vm_group_bin_15495 = frame (4k)
frame_vm_group_bin_15496 = frame (4k)
frame_vm_group_bin_15497 = frame (4k)
frame_vm_group_bin_15498 = frame (4k)
frame_vm_group_bin_15499 = frame (4k)
frame_vm_group_bin_1550 = frame (4k)
frame_vm_group_bin_15500 = frame (4k)
frame_vm_group_bin_15501 = frame (4k)
frame_vm_group_bin_15502 = frame (4k)
frame_vm_group_bin_15503 = frame (4k)
frame_vm_group_bin_15504 = frame (4k)
frame_vm_group_bin_15505 = frame (4k)
frame_vm_group_bin_15506 = frame (4k)
frame_vm_group_bin_15507 = frame (4k)
frame_vm_group_bin_15508 = frame (4k)
frame_vm_group_bin_15509 = frame (4k)
frame_vm_group_bin_1551 = frame (4k)
frame_vm_group_bin_15510 = frame (4k)
frame_vm_group_bin_15511 = frame (4k)
frame_vm_group_bin_15512 = frame (4k)
frame_vm_group_bin_15513 = frame (4k)
frame_vm_group_bin_15514 = frame (4k)
frame_vm_group_bin_15515 = frame (4k)
frame_vm_group_bin_15516 = frame (4k)
frame_vm_group_bin_15517 = frame (4k)
frame_vm_group_bin_15518 = frame (4k)
frame_vm_group_bin_15519 = frame (4k)
frame_vm_group_bin_1552 = frame (4k)
frame_vm_group_bin_15520 = frame (4k)
frame_vm_group_bin_15521 = frame (4k)
frame_vm_group_bin_15522 = frame (4k)
frame_vm_group_bin_15523 = frame (4k)
frame_vm_group_bin_15524 = frame (4k)
frame_vm_group_bin_15525 = frame (4k)
frame_vm_group_bin_15526 = frame (4k)
frame_vm_group_bin_15527 = frame (4k)
frame_vm_group_bin_15528 = frame (4k)
frame_vm_group_bin_15529 = frame (4k)
frame_vm_group_bin_1553 = frame (4k)
frame_vm_group_bin_15530 = frame (4k)
frame_vm_group_bin_15531 = frame (4k)
frame_vm_group_bin_15532 = frame (4k)
frame_vm_group_bin_15533 = frame (4k)
frame_vm_group_bin_15534 = frame (4k)
frame_vm_group_bin_15535 = frame (4k)
frame_vm_group_bin_15536 = frame (4k)
frame_vm_group_bin_15537 = frame (4k)
frame_vm_group_bin_15538 = frame (4k)
frame_vm_group_bin_15539 = frame (4k)
frame_vm_group_bin_1554 = frame (4k)
frame_vm_group_bin_15540 = frame (4k)
frame_vm_group_bin_15541 = frame (4k)
frame_vm_group_bin_15542 = frame (4k)
frame_vm_group_bin_15543 = frame (4k)
frame_vm_group_bin_15544 = frame (4k)
frame_vm_group_bin_15545 = frame (4k)
frame_vm_group_bin_15546 = frame (4k)
frame_vm_group_bin_15547 = frame (4k)
frame_vm_group_bin_15548 = frame (4k)
frame_vm_group_bin_15549 = frame (4k)
frame_vm_group_bin_1555 = frame (4k)
frame_vm_group_bin_15550 = frame (4k)
frame_vm_group_bin_15551 = frame (4k)
frame_vm_group_bin_15552 = frame (4k)
frame_vm_group_bin_15553 = frame (4k)
frame_vm_group_bin_15554 = frame (4k)
frame_vm_group_bin_15555 = frame (4k)
frame_vm_group_bin_15556 = frame (4k)
frame_vm_group_bin_15557 = frame (4k)
frame_vm_group_bin_15558 = frame (4k)
frame_vm_group_bin_15559 = frame (4k)
frame_vm_group_bin_1556 = frame (4k)
frame_vm_group_bin_15560 = frame (4k)
frame_vm_group_bin_15561 = frame (4k)
frame_vm_group_bin_15562 = frame (4k)
frame_vm_group_bin_15563 = frame (4k)
frame_vm_group_bin_15564 = frame (4k)
frame_vm_group_bin_15565 = frame (4k)
frame_vm_group_bin_15566 = frame (4k)
frame_vm_group_bin_15567 = frame (4k)
frame_vm_group_bin_15568 = frame (4k)
frame_vm_group_bin_15569 = frame (4k)
frame_vm_group_bin_1557 = frame (4k)
frame_vm_group_bin_15570 = frame (4k)
frame_vm_group_bin_15571 = frame (4k)
frame_vm_group_bin_15572 = frame (4k)
frame_vm_group_bin_15573 = frame (4k)
frame_vm_group_bin_15574 = frame (4k)
frame_vm_group_bin_15575 = frame (4k)
frame_vm_group_bin_15576 = frame (4k)
frame_vm_group_bin_15577 = frame (4k)
frame_vm_group_bin_15578 = frame (4k)
frame_vm_group_bin_15579 = frame (4k)
frame_vm_group_bin_1558 = frame (4k)
frame_vm_group_bin_15580 = frame (4k)
frame_vm_group_bin_15581 = frame (4k)
frame_vm_group_bin_15582 = frame (4k)
frame_vm_group_bin_15583 = frame (4k)
frame_vm_group_bin_15584 = frame (4k)
frame_vm_group_bin_15585 = frame (4k)
frame_vm_group_bin_15586 = frame (4k)
frame_vm_group_bin_15587 = frame (4k)
frame_vm_group_bin_15588 = frame (4k)
frame_vm_group_bin_15589 = frame (4k)
frame_vm_group_bin_1559 = frame (4k)
frame_vm_group_bin_15590 = frame (4k)
frame_vm_group_bin_15591 = frame (4k)
frame_vm_group_bin_15592 = frame (4k)
frame_vm_group_bin_15593 = frame (4k)
frame_vm_group_bin_15594 = frame (4k)
frame_vm_group_bin_15595 = frame (4k)
frame_vm_group_bin_15596 = frame (4k)
frame_vm_group_bin_15597 = frame (4k)
frame_vm_group_bin_15598 = frame (4k)
frame_vm_group_bin_15599 = frame (4k)
frame_vm_group_bin_1560 = frame (4k)
frame_vm_group_bin_15600 = frame (4k)
frame_vm_group_bin_15601 = frame (4k)
frame_vm_group_bin_15602 = frame (4k)
frame_vm_group_bin_15603 = frame (4k)
frame_vm_group_bin_15604 = frame (4k)
frame_vm_group_bin_15605 = frame (4k)
frame_vm_group_bin_15606 = frame (4k)
frame_vm_group_bin_15607 = frame (4k)
frame_vm_group_bin_15608 = frame (4k)
frame_vm_group_bin_15609 = frame (4k)
frame_vm_group_bin_1561 = frame (4k)
frame_vm_group_bin_15610 = frame (4k)
frame_vm_group_bin_15611 = frame (4k)
frame_vm_group_bin_15612 = frame (4k)
frame_vm_group_bin_15613 = frame (4k)
frame_vm_group_bin_15614 = frame (4k)
frame_vm_group_bin_15615 = frame (4k)
frame_vm_group_bin_15616 = frame (4k)
frame_vm_group_bin_15617 = frame (4k)
frame_vm_group_bin_15618 = frame (4k)
frame_vm_group_bin_15619 = frame (4k)
frame_vm_group_bin_1562 = frame (4k)
frame_vm_group_bin_15620 = frame (4k)
frame_vm_group_bin_15621 = frame (4k)
frame_vm_group_bin_15622 = frame (4k)
frame_vm_group_bin_15623 = frame (4k)
frame_vm_group_bin_15624 = frame (4k)
frame_vm_group_bin_15625 = frame (4k)
frame_vm_group_bin_15626 = frame (4k)
frame_vm_group_bin_15627 = frame (4k)
frame_vm_group_bin_15628 = frame (4k)
frame_vm_group_bin_15629 = frame (4k)
frame_vm_group_bin_1563 = frame (4k)
frame_vm_group_bin_15630 = frame (4k)
frame_vm_group_bin_15631 = frame (4k)
frame_vm_group_bin_15632 = frame (4k)
frame_vm_group_bin_15633 = frame (4k)
frame_vm_group_bin_15634 = frame (4k)
frame_vm_group_bin_15635 = frame (4k)
frame_vm_group_bin_15636 = frame (4k)
frame_vm_group_bin_15637 = frame (4k)
frame_vm_group_bin_15638 = frame (4k)
frame_vm_group_bin_15639 = frame (4k)
frame_vm_group_bin_1564 = frame (4k)
frame_vm_group_bin_15640 = frame (4k)
frame_vm_group_bin_15641 = frame (4k)
frame_vm_group_bin_15642 = frame (4k)
frame_vm_group_bin_15643 = frame (4k)
frame_vm_group_bin_15644 = frame (4k)
frame_vm_group_bin_15645 = frame (4k)
frame_vm_group_bin_15646 = frame (4k)
frame_vm_group_bin_15647 = frame (4k)
frame_vm_group_bin_15648 = frame (4k)
frame_vm_group_bin_15649 = frame (4k)
frame_vm_group_bin_1565 = frame (4k)
frame_vm_group_bin_15650 = frame (4k)
frame_vm_group_bin_15651 = frame (4k)
frame_vm_group_bin_15652 = frame (4k)
frame_vm_group_bin_15653 = frame (4k)
frame_vm_group_bin_15654 = frame (4k)
frame_vm_group_bin_15655 = frame (4k)
frame_vm_group_bin_15656 = frame (4k)
frame_vm_group_bin_15657 = frame (4k)
frame_vm_group_bin_15658 = frame (4k)
frame_vm_group_bin_15659 = frame (4k)
frame_vm_group_bin_1566 = frame (4k)
frame_vm_group_bin_15660 = frame (4k)
frame_vm_group_bin_15661 = frame (4k)
frame_vm_group_bin_15662 = frame (4k)
frame_vm_group_bin_15663 = frame (4k)
frame_vm_group_bin_15664 = frame (4k)
frame_vm_group_bin_15665 = frame (4k)
frame_vm_group_bin_15666 = frame (4k)
frame_vm_group_bin_15667 = frame (4k)
frame_vm_group_bin_15668 = frame (4k)
frame_vm_group_bin_15669 = frame (4k)
frame_vm_group_bin_1567 = frame (4k)
frame_vm_group_bin_15670 = frame (4k)
frame_vm_group_bin_15671 = frame (4k)
frame_vm_group_bin_15672 = frame (4k)
frame_vm_group_bin_15673 = frame (4k)
frame_vm_group_bin_15674 = frame (4k)
frame_vm_group_bin_15675 = frame (4k)
frame_vm_group_bin_15676 = frame (4k)
frame_vm_group_bin_15677 = frame (4k)
frame_vm_group_bin_15678 = frame (4k)
frame_vm_group_bin_15679 = frame (4k)
frame_vm_group_bin_1568 = frame (4k)
frame_vm_group_bin_15680 = frame (4k)
frame_vm_group_bin_15681 = frame (4k)
frame_vm_group_bin_15682 = frame (4k)
frame_vm_group_bin_15683 = frame (4k)
frame_vm_group_bin_15684 = frame (4k)
frame_vm_group_bin_15685 = frame (4k)
frame_vm_group_bin_15686 = frame (4k)
frame_vm_group_bin_15687 = frame (4k)
frame_vm_group_bin_15688 = frame (4k)
frame_vm_group_bin_15689 = frame (4k)
frame_vm_group_bin_1569 = frame (4k)
frame_vm_group_bin_15690 = frame (4k)
frame_vm_group_bin_15691 = frame (4k)
frame_vm_group_bin_15692 = frame (4k)
frame_vm_group_bin_15693 = frame (4k)
frame_vm_group_bin_15694 = frame (4k)
frame_vm_group_bin_15695 = frame (4k)
frame_vm_group_bin_15696 = frame (4k)
frame_vm_group_bin_15697 = frame (4k)
frame_vm_group_bin_15698 = frame (4k)
frame_vm_group_bin_15699 = frame (4k)
frame_vm_group_bin_1570 = frame (4k)
frame_vm_group_bin_15700 = frame (4k)
frame_vm_group_bin_15701 = frame (4k)
frame_vm_group_bin_15702 = frame (4k)
frame_vm_group_bin_15703 = frame (4k)
frame_vm_group_bin_15704 = frame (4k)
frame_vm_group_bin_15705 = frame (4k)
frame_vm_group_bin_15706 = frame (4k)
frame_vm_group_bin_15707 = frame (4k)
frame_vm_group_bin_15708 = frame (4k)
frame_vm_group_bin_15709 = frame (4k)
frame_vm_group_bin_1571 = frame (4k)
frame_vm_group_bin_15710 = frame (4k)
frame_vm_group_bin_15711 = frame (4k)
frame_vm_group_bin_15712 = frame (4k)
frame_vm_group_bin_15713 = frame (4k)
frame_vm_group_bin_15714 = frame (4k)
frame_vm_group_bin_15715 = frame (4k)
frame_vm_group_bin_15716 = frame (4k)
frame_vm_group_bin_15717 = frame (4k)
frame_vm_group_bin_15718 = frame (4k)
frame_vm_group_bin_15719 = frame (4k)
frame_vm_group_bin_1572 = frame (4k)
frame_vm_group_bin_15720 = frame (4k)
frame_vm_group_bin_15721 = frame (4k)
frame_vm_group_bin_15722 = frame (4k)
frame_vm_group_bin_15723 = frame (4k)
frame_vm_group_bin_15724 = frame (4k)
frame_vm_group_bin_15725 = frame (4k)
frame_vm_group_bin_15726 = frame (4k)
frame_vm_group_bin_15727 = frame (4k)
frame_vm_group_bin_15728 = frame (4k)
frame_vm_group_bin_15729 = frame (4k)
frame_vm_group_bin_1573 = frame (4k)
frame_vm_group_bin_15730 = frame (4k)
frame_vm_group_bin_15731 = frame (4k)
frame_vm_group_bin_15732 = frame (4k)
frame_vm_group_bin_15733 = frame (4k)
frame_vm_group_bin_15734 = frame (4k)
frame_vm_group_bin_15735 = frame (4k)
frame_vm_group_bin_15736 = frame (4k)
frame_vm_group_bin_15737 = frame (4k)
frame_vm_group_bin_15738 = frame (4k)
frame_vm_group_bin_15739 = frame (4k)
frame_vm_group_bin_1574 = frame (4k)
frame_vm_group_bin_15740 = frame (4k)
frame_vm_group_bin_15741 = frame (4k)
frame_vm_group_bin_15742 = frame (4k)
frame_vm_group_bin_15743 = frame (4k)
frame_vm_group_bin_15744 = frame (4k)
frame_vm_group_bin_15745 = frame (4k)
frame_vm_group_bin_15746 = frame (4k)
frame_vm_group_bin_15747 = frame (4k)
frame_vm_group_bin_15748 = frame (4k)
frame_vm_group_bin_15749 = frame (4k)
frame_vm_group_bin_1575 = frame (4k)
frame_vm_group_bin_15750 = frame (4k)
frame_vm_group_bin_15751 = frame (4k)
frame_vm_group_bin_15752 = frame (4k)
frame_vm_group_bin_15753 = frame (4k)
frame_vm_group_bin_15754 = frame (4k)
frame_vm_group_bin_15755 = frame (4k)
frame_vm_group_bin_15756 = frame (4k)
frame_vm_group_bin_15757 = frame (4k)
frame_vm_group_bin_15758 = frame (4k)
frame_vm_group_bin_15759 = frame (4k)
frame_vm_group_bin_1576 = frame (4k)
frame_vm_group_bin_15760 = frame (4k)
frame_vm_group_bin_15761 = frame (4k)
frame_vm_group_bin_15762 = frame (4k)
frame_vm_group_bin_15763 = frame (4k)
frame_vm_group_bin_15764 = frame (4k)
frame_vm_group_bin_15765 = frame (4k)
frame_vm_group_bin_15766 = frame (4k)
frame_vm_group_bin_15767 = frame (4k)
frame_vm_group_bin_15768 = frame (4k)
frame_vm_group_bin_15769 = frame (4k)
frame_vm_group_bin_1577 = frame (4k)
frame_vm_group_bin_15770 = frame (4k)
frame_vm_group_bin_15771 = frame (4k)
frame_vm_group_bin_15772 = frame (4k)
frame_vm_group_bin_15773 = frame (4k)
frame_vm_group_bin_15774 = frame (4k)
frame_vm_group_bin_15775 = frame (4k)
frame_vm_group_bin_15776 = frame (4k)
frame_vm_group_bin_15777 = frame (4k)
frame_vm_group_bin_15778 = frame (4k)
frame_vm_group_bin_15779 = frame (4k)
frame_vm_group_bin_1578 = frame (4k)
frame_vm_group_bin_15780 = frame (4k)
frame_vm_group_bin_15781 = frame (4k)
frame_vm_group_bin_15782 = frame (4k)
frame_vm_group_bin_15783 = frame (4k)
frame_vm_group_bin_15784 = frame (4k)
frame_vm_group_bin_15785 = frame (4k)
frame_vm_group_bin_15786 = frame (4k)
frame_vm_group_bin_15787 = frame (4k)
frame_vm_group_bin_15788 = frame (4k)
frame_vm_group_bin_15789 = frame (4k)
frame_vm_group_bin_1579 = frame (4k)
frame_vm_group_bin_15790 = frame (4k)
frame_vm_group_bin_15791 = frame (4k)
frame_vm_group_bin_15792 = frame (4k)
frame_vm_group_bin_15793 = frame (4k)
frame_vm_group_bin_15794 = frame (4k)
frame_vm_group_bin_15795 = frame (4k)
frame_vm_group_bin_15796 = frame (4k)
frame_vm_group_bin_15797 = frame (4k)
frame_vm_group_bin_15798 = frame (4k)
frame_vm_group_bin_15799 = frame (4k)
frame_vm_group_bin_1580 = frame (4k)
frame_vm_group_bin_15800 = frame (4k)
frame_vm_group_bin_15801 = frame (4k)
frame_vm_group_bin_15802 = frame (4k)
frame_vm_group_bin_15803 = frame (4k)
frame_vm_group_bin_15804 = frame (4k)
frame_vm_group_bin_15805 = frame (4k)
frame_vm_group_bin_15806 = frame (4k)
frame_vm_group_bin_15807 = frame (4k)
frame_vm_group_bin_15808 = frame (4k)
frame_vm_group_bin_15809 = frame (4k)
frame_vm_group_bin_1581 = frame (4k)
frame_vm_group_bin_15810 = frame (4k)
frame_vm_group_bin_15811 = frame (4k)
frame_vm_group_bin_15812 = frame (4k)
frame_vm_group_bin_15813 = frame (4k)
frame_vm_group_bin_15814 = frame (4k)
frame_vm_group_bin_15815 = frame (4k)
frame_vm_group_bin_15816 = frame (4k)
frame_vm_group_bin_15817 = frame (4k)
frame_vm_group_bin_15818 = frame (4k)
frame_vm_group_bin_15819 = frame (4k)
frame_vm_group_bin_1582 = frame (4k)
frame_vm_group_bin_15820 = frame (4k)
frame_vm_group_bin_15821 = frame (4k)
frame_vm_group_bin_15822 = frame (4k)
frame_vm_group_bin_15823 = frame (4k)
frame_vm_group_bin_15824 = frame (4k)
frame_vm_group_bin_15825 = frame (4k)
frame_vm_group_bin_15826 = frame (4k)
frame_vm_group_bin_15827 = frame (4k)
frame_vm_group_bin_15828 = frame (4k)
frame_vm_group_bin_15829 = frame (4k)
frame_vm_group_bin_1583 = frame (4k)
frame_vm_group_bin_15830 = frame (4k)
frame_vm_group_bin_15831 = frame (4k)
frame_vm_group_bin_15832 = frame (4k)
frame_vm_group_bin_15833 = frame (4k)
frame_vm_group_bin_15834 = frame (4k)
frame_vm_group_bin_15835 = frame (4k)
frame_vm_group_bin_15836 = frame (4k)
frame_vm_group_bin_15837 = frame (4k)
frame_vm_group_bin_15838 = frame (4k)
frame_vm_group_bin_15839 = frame (4k)
frame_vm_group_bin_1584 = frame (4k)
frame_vm_group_bin_15840 = frame (4k)
frame_vm_group_bin_15841 = frame (4k)
frame_vm_group_bin_15842 = frame (4k)
frame_vm_group_bin_15843 = frame (4k)
frame_vm_group_bin_15844 = frame (4k)
frame_vm_group_bin_15845 = frame (4k)
frame_vm_group_bin_15846 = frame (4k)
frame_vm_group_bin_15847 = frame (4k)
frame_vm_group_bin_15848 = frame (4k)
frame_vm_group_bin_15849 = frame (4k)
frame_vm_group_bin_1585 = frame (4k)
frame_vm_group_bin_15850 = frame (4k)
frame_vm_group_bin_15851 = frame (4k)
frame_vm_group_bin_15852 = frame (4k)
frame_vm_group_bin_15853 = frame (4k)
frame_vm_group_bin_15854 = frame (4k)
frame_vm_group_bin_15855 = frame (4k)
frame_vm_group_bin_15856 = frame (4k)
frame_vm_group_bin_15857 = frame (4k)
frame_vm_group_bin_15858 = frame (4k)
frame_vm_group_bin_15859 = frame (4k)
frame_vm_group_bin_1586 = frame (4k)
frame_vm_group_bin_15860 = frame (4k)
frame_vm_group_bin_15861 = frame (4k)
frame_vm_group_bin_15862 = frame (4k)
frame_vm_group_bin_15863 = frame (4k)
frame_vm_group_bin_15864 = frame (4k)
frame_vm_group_bin_15865 = frame (4k)
frame_vm_group_bin_15866 = frame (4k)
frame_vm_group_bin_15867 = frame (4k)
frame_vm_group_bin_15868 = frame (4k)
frame_vm_group_bin_15869 = frame (4k)
frame_vm_group_bin_1587 = frame (4k)
frame_vm_group_bin_15870 = frame (4k)
frame_vm_group_bin_15871 = frame (4k)
frame_vm_group_bin_15872 = frame (4k)
frame_vm_group_bin_15873 = frame (4k)
frame_vm_group_bin_15874 = frame (4k)
frame_vm_group_bin_15875 = frame (4k)
frame_vm_group_bin_15876 = frame (4k)
frame_vm_group_bin_15877 = frame (4k)
frame_vm_group_bin_15878 = frame (4k)
frame_vm_group_bin_15879 = frame (4k)
frame_vm_group_bin_1588 = frame (4k)
frame_vm_group_bin_15880 = frame (4k)
frame_vm_group_bin_15881 = frame (4k)
frame_vm_group_bin_15882 = frame (4k)
frame_vm_group_bin_15883 = frame (4k)
frame_vm_group_bin_15884 = frame (4k)
frame_vm_group_bin_15885 = frame (4k)
frame_vm_group_bin_15886 = frame (4k)
frame_vm_group_bin_15887 = frame (4k)
frame_vm_group_bin_15888 = frame (4k)
frame_vm_group_bin_15889 = frame (4k)
frame_vm_group_bin_1589 = frame (4k)
frame_vm_group_bin_15890 = frame (4k)
frame_vm_group_bin_15891 = frame (4k)
frame_vm_group_bin_15892 = frame (4k)
frame_vm_group_bin_15893 = frame (4k)
frame_vm_group_bin_15894 = frame (4k)
frame_vm_group_bin_15895 = frame (4k)
frame_vm_group_bin_15896 = frame (4k)
frame_vm_group_bin_15897 = frame (4k)
frame_vm_group_bin_15898 = frame (4k)
frame_vm_group_bin_15899 = frame (4k)
frame_vm_group_bin_1590 = frame (4k)
frame_vm_group_bin_15900 = frame (4k)
frame_vm_group_bin_15901 = frame (4k)
frame_vm_group_bin_15902 = frame (4k)
frame_vm_group_bin_15903 = frame (4k)
frame_vm_group_bin_15904 = frame (4k)
frame_vm_group_bin_15905 = frame (4k)
frame_vm_group_bin_15906 = frame (4k)
frame_vm_group_bin_15907 = frame (4k)
frame_vm_group_bin_15908 = frame (4k)
frame_vm_group_bin_15909 = frame (4k)
frame_vm_group_bin_1591 = frame (4k)
frame_vm_group_bin_15910 = frame (4k)
frame_vm_group_bin_15911 = frame (4k)
frame_vm_group_bin_15912 = frame (4k)
frame_vm_group_bin_15913 = frame (4k)
frame_vm_group_bin_15914 = frame (4k)
frame_vm_group_bin_15915 = frame (4k)
frame_vm_group_bin_15916 = frame (4k)
frame_vm_group_bin_15917 = frame (4k)
frame_vm_group_bin_15918 = frame (4k)
frame_vm_group_bin_15919 = frame (4k)
frame_vm_group_bin_1592 = frame (4k)
frame_vm_group_bin_15920 = frame (4k)
frame_vm_group_bin_15921 = frame (4k)
frame_vm_group_bin_15922 = frame (4k)
frame_vm_group_bin_15923 = frame (4k)
frame_vm_group_bin_15924 = frame (4k)
frame_vm_group_bin_15925 = frame (4k)
frame_vm_group_bin_15926 = frame (4k)
frame_vm_group_bin_15927 = frame (4k)
frame_vm_group_bin_15928 = frame (4k)
frame_vm_group_bin_15929 = frame (4k)
frame_vm_group_bin_1593 = frame (4k)
frame_vm_group_bin_15930 = frame (4k)
frame_vm_group_bin_15931 = frame (4k)
frame_vm_group_bin_15932 = frame (4k)
frame_vm_group_bin_15933 = frame (4k)
frame_vm_group_bin_15934 = frame (4k)
frame_vm_group_bin_15935 = frame (4k)
frame_vm_group_bin_15936 = frame (4k)
frame_vm_group_bin_15937 = frame (4k)
frame_vm_group_bin_15938 = frame (4k)
frame_vm_group_bin_15939 = frame (4k)
frame_vm_group_bin_1594 = frame (4k)
frame_vm_group_bin_15940 = frame (4k)
frame_vm_group_bin_15941 = frame (4k)
frame_vm_group_bin_15942 = frame (4k)
frame_vm_group_bin_15943 = frame (4k)
frame_vm_group_bin_15944 = frame (4k)
frame_vm_group_bin_15945 = frame (4k)
frame_vm_group_bin_15946 = frame (4k)
frame_vm_group_bin_15947 = frame (4k)
frame_vm_group_bin_15948 = frame (4k)
frame_vm_group_bin_15949 = frame (4k)
frame_vm_group_bin_1595 = frame (4k)
frame_vm_group_bin_15950 = frame (4k)
frame_vm_group_bin_15951 = frame (4k)
frame_vm_group_bin_15952 = frame (4k)
frame_vm_group_bin_15953 = frame (4k)
frame_vm_group_bin_15954 = frame (4k)
frame_vm_group_bin_15955 = frame (4k)
frame_vm_group_bin_15956 = frame (4k)
frame_vm_group_bin_15957 = frame (4k)
frame_vm_group_bin_15958 = frame (4k)
frame_vm_group_bin_15959 = frame (4k)
frame_vm_group_bin_1596 = frame (4k)
frame_vm_group_bin_15960 = frame (4k)
frame_vm_group_bin_15961 = frame (4k)
frame_vm_group_bin_15962 = frame (4k)
frame_vm_group_bin_15963 = frame (4k)
frame_vm_group_bin_15964 = frame (4k)
frame_vm_group_bin_15965 = frame (4k)
frame_vm_group_bin_15966 = frame (4k)
frame_vm_group_bin_15967 = frame (4k)
frame_vm_group_bin_15968 = frame (4k)
frame_vm_group_bin_15969 = frame (4k)
frame_vm_group_bin_1597 = frame (4k)
frame_vm_group_bin_15970 = frame (4k)
frame_vm_group_bin_15971 = frame (4k)
frame_vm_group_bin_15972 = frame (4k)
frame_vm_group_bin_15973 = frame (4k)
frame_vm_group_bin_15974 = frame (4k)
frame_vm_group_bin_15975 = frame (4k)
frame_vm_group_bin_15976 = frame (4k)
frame_vm_group_bin_15977 = frame (4k)
frame_vm_group_bin_15978 = frame (4k)
frame_vm_group_bin_15979 = frame (4k)
frame_vm_group_bin_1598 = frame (4k)
frame_vm_group_bin_15980 = frame (4k)
frame_vm_group_bin_15981 = frame (4k)
frame_vm_group_bin_15982 = frame (4k)
frame_vm_group_bin_15983 = frame (4k)
frame_vm_group_bin_15984 = frame (4k)
frame_vm_group_bin_15985 = frame (4k)
frame_vm_group_bin_15986 = frame (4k)
frame_vm_group_bin_15987 = frame (4k)
frame_vm_group_bin_15988 = frame (4k)
frame_vm_group_bin_15989 = frame (4k)
frame_vm_group_bin_1599 = frame (4k)
frame_vm_group_bin_15990 = frame (4k)
frame_vm_group_bin_15991 = frame (4k)
frame_vm_group_bin_15992 = frame (4k)
frame_vm_group_bin_15993 = frame (4k)
frame_vm_group_bin_15994 = frame (4k)
frame_vm_group_bin_15995 = frame (4k)
frame_vm_group_bin_15996 = frame (4k)
frame_vm_group_bin_15997 = frame (4k)
frame_vm_group_bin_15998 = frame (4k)
frame_vm_group_bin_15999 = frame (4k)
frame_vm_group_bin_1600 = frame (4k)
frame_vm_group_bin_16000 = frame (4k)
frame_vm_group_bin_16001 = frame (4k)
frame_vm_group_bin_16002 = frame (4k)
frame_vm_group_bin_16003 = frame (4k)
frame_vm_group_bin_16004 = frame (4k)
frame_vm_group_bin_16005 = frame (4k)
frame_vm_group_bin_16006 = frame (4k)
frame_vm_group_bin_16007 = frame (4k)
frame_vm_group_bin_16008 = frame (4k)
frame_vm_group_bin_16009 = frame (4k)
frame_vm_group_bin_1601 = frame (4k)
frame_vm_group_bin_16010 = frame (4k)
frame_vm_group_bin_16011 = frame (4k)
frame_vm_group_bin_16012 = frame (4k)
frame_vm_group_bin_16013 = frame (4k)
frame_vm_group_bin_16014 = frame (4k)
frame_vm_group_bin_16016 = frame (4k)
frame_vm_group_bin_16017 = frame (4k)
frame_vm_group_bin_16018 = frame (4k)
frame_vm_group_bin_16019 = frame (4k)
frame_vm_group_bin_1602 = frame (4k)
frame_vm_group_bin_16020 = frame (4k)
frame_vm_group_bin_16021 = frame (4k)
frame_vm_group_bin_16022 = frame (4k)
frame_vm_group_bin_16023 = frame (4k)
frame_vm_group_bin_16024 = frame (4k)
frame_vm_group_bin_16025 = frame (4k)
frame_vm_group_bin_16026 = frame (4k)
frame_vm_group_bin_16027 = frame (4k)
frame_vm_group_bin_16028 = frame (4k)
frame_vm_group_bin_16029 = frame (4k)
frame_vm_group_bin_1603 = frame (4k)
frame_vm_group_bin_16030 = frame (4k)
frame_vm_group_bin_16031 = frame (4k)
frame_vm_group_bin_16032 = frame (4k)
frame_vm_group_bin_16033 = frame (4k)
frame_vm_group_bin_16034 = frame (4k)
frame_vm_group_bin_16035 = frame (4k)
frame_vm_group_bin_16036 = frame (4k)
frame_vm_group_bin_16037 = frame (4k)
frame_vm_group_bin_16038 = frame (4k)
frame_vm_group_bin_16039 = frame (4k)
frame_vm_group_bin_1604 = frame (4k)
frame_vm_group_bin_16040 = frame (4k)
frame_vm_group_bin_16041 = frame (4k)
frame_vm_group_bin_16042 = frame (4k)
frame_vm_group_bin_16043 = frame (4k)
frame_vm_group_bin_16044 = frame (4k)
frame_vm_group_bin_16045 = frame (4k)
frame_vm_group_bin_16046 = frame (4k)
frame_vm_group_bin_16047 = frame (4k)
frame_vm_group_bin_16048 = frame (4k)
frame_vm_group_bin_16049 = frame (4k)
frame_vm_group_bin_1605 = frame (4k)
frame_vm_group_bin_16050 = frame (4k)
frame_vm_group_bin_16051 = frame (4k)
frame_vm_group_bin_16052 = frame (4k)
frame_vm_group_bin_16053 = frame (4k)
frame_vm_group_bin_16054 = frame (4k)
frame_vm_group_bin_16055 = frame (4k)
frame_vm_group_bin_16056 = frame (4k)
frame_vm_group_bin_16057 = frame (4k)
frame_vm_group_bin_16058 = frame (4k)
frame_vm_group_bin_16059 = frame (4k)
frame_vm_group_bin_1606 = frame (4k)
frame_vm_group_bin_16060 = frame (4k)
frame_vm_group_bin_16061 = frame (4k)
frame_vm_group_bin_16062 = frame (4k)
frame_vm_group_bin_16063 = frame (4k)
frame_vm_group_bin_16064 = frame (4k)
frame_vm_group_bin_16065 = frame (4k)
frame_vm_group_bin_16066 = frame (4k)
frame_vm_group_bin_16067 = frame (4k)
frame_vm_group_bin_16068 = frame (4k)
frame_vm_group_bin_16069 = frame (4k)
frame_vm_group_bin_1607 = frame (4k)
frame_vm_group_bin_16070 = frame (4k)
frame_vm_group_bin_16071 = frame (4k)
frame_vm_group_bin_16072 = frame (4k)
frame_vm_group_bin_16073 = frame (4k)
frame_vm_group_bin_16074 = frame (4k)
frame_vm_group_bin_16075 = frame (4k)
frame_vm_group_bin_16076 = frame (4k)
frame_vm_group_bin_16077 = frame (4k)
frame_vm_group_bin_16078 = frame (4k)
frame_vm_group_bin_16079 = frame (4k)
frame_vm_group_bin_1608 = frame (4k)
frame_vm_group_bin_16080 = frame (4k)
frame_vm_group_bin_16081 = frame (4k)
frame_vm_group_bin_16082 = frame (4k)
frame_vm_group_bin_16083 = frame (4k)
frame_vm_group_bin_16084 = frame (4k)
frame_vm_group_bin_16085 = frame (4k)
frame_vm_group_bin_16086 = frame (4k)
frame_vm_group_bin_16087 = frame (4k)
frame_vm_group_bin_16088 = frame (4k)
frame_vm_group_bin_16089 = frame (4k)
frame_vm_group_bin_1609 = frame (4k)
frame_vm_group_bin_16090 = frame (4k)
frame_vm_group_bin_16091 = frame (4k)
frame_vm_group_bin_16092 = frame (4k)
frame_vm_group_bin_16093 = frame (4k)
frame_vm_group_bin_16094 = frame (4k)
frame_vm_group_bin_16095 = frame (4k)
frame_vm_group_bin_16096 = frame (4k)
frame_vm_group_bin_16097 = frame (4k)
frame_vm_group_bin_16098 = frame (4k)
frame_vm_group_bin_16099 = frame (4k)
frame_vm_group_bin_1610 = frame (4k)
frame_vm_group_bin_16100 = frame (4k)
frame_vm_group_bin_16101 = frame (4k)
frame_vm_group_bin_16102 = frame (4k)
frame_vm_group_bin_16103 = frame (4k)
frame_vm_group_bin_16104 = frame (4k)
frame_vm_group_bin_16105 = frame (4k)
frame_vm_group_bin_16106 = frame (4k)
frame_vm_group_bin_16107 = frame (4k)
frame_vm_group_bin_16108 = frame (4k)
frame_vm_group_bin_16109 = frame (4k)
frame_vm_group_bin_1611 = frame (4k)
frame_vm_group_bin_16110 = frame (4k)
frame_vm_group_bin_16111 = frame (4k)
frame_vm_group_bin_16112 = frame (4k)
frame_vm_group_bin_16113 = frame (4k)
frame_vm_group_bin_16114 = frame (4k)
frame_vm_group_bin_16115 = frame (4k)
frame_vm_group_bin_16116 = frame (4k)
frame_vm_group_bin_16117 = frame (4k)
frame_vm_group_bin_16118 = frame (4k)
frame_vm_group_bin_16119 = frame (4k)
frame_vm_group_bin_1612 = frame (4k)
frame_vm_group_bin_16120 = frame (4k)
frame_vm_group_bin_16121 = frame (4k)
frame_vm_group_bin_16122 = frame (4k)
frame_vm_group_bin_16123 = frame (4k)
frame_vm_group_bin_16124 = frame (4k)
frame_vm_group_bin_16125 = frame (4k)
frame_vm_group_bin_16126 = frame (4k)
frame_vm_group_bin_16127 = frame (4k)
frame_vm_group_bin_16128 = frame (4k)
frame_vm_group_bin_16129 = frame (4k)
frame_vm_group_bin_1613 = frame (4k)
frame_vm_group_bin_16130 = frame (4k)
frame_vm_group_bin_16131 = frame (4k)
frame_vm_group_bin_16132 = frame (4k)
frame_vm_group_bin_16133 = frame (4k)
frame_vm_group_bin_16134 = frame (4k)
frame_vm_group_bin_16135 = frame (4k)
frame_vm_group_bin_16136 = frame (4k)
frame_vm_group_bin_16137 = frame (4k)
frame_vm_group_bin_16138 = frame (4k)
frame_vm_group_bin_16139 = frame (4k)
frame_vm_group_bin_1614 = frame (4k)
frame_vm_group_bin_16140 = frame (4k)
frame_vm_group_bin_16141 = frame (4k)
frame_vm_group_bin_16142 = frame (4k)
frame_vm_group_bin_16143 = frame (4k)
frame_vm_group_bin_16144 = frame (4k)
frame_vm_group_bin_16145 = frame (4k)
frame_vm_group_bin_16146 = frame (4k)
frame_vm_group_bin_16147 = frame (4k)
frame_vm_group_bin_16148 = frame (4k)
frame_vm_group_bin_16149 = frame (4k)
frame_vm_group_bin_1615 = frame (4k)
frame_vm_group_bin_16150 = frame (4k)
frame_vm_group_bin_16151 = frame (4k)
frame_vm_group_bin_16152 = frame (4k)
frame_vm_group_bin_16153 = frame (4k)
frame_vm_group_bin_16154 = frame (4k)
frame_vm_group_bin_16155 = frame (4k)
frame_vm_group_bin_16156 = frame (4k)
frame_vm_group_bin_16157 = frame (4k)
frame_vm_group_bin_16158 = frame (4k)
frame_vm_group_bin_16159 = frame (4k)
frame_vm_group_bin_1616 = frame (4k)
frame_vm_group_bin_16160 = frame (4k)
frame_vm_group_bin_16161 = frame (4k)
frame_vm_group_bin_16162 = frame (4k)
frame_vm_group_bin_16163 = frame (4k)
frame_vm_group_bin_16164 = frame (4k)
frame_vm_group_bin_16165 = frame (4k)
frame_vm_group_bin_16166 = frame (4k)
frame_vm_group_bin_16167 = frame (4k)
frame_vm_group_bin_16168 = frame (4k)
frame_vm_group_bin_16169 = frame (4k)
frame_vm_group_bin_1617 = frame (4k)
frame_vm_group_bin_16170 = frame (4k)
frame_vm_group_bin_16171 = frame (4k)
frame_vm_group_bin_16172 = frame (4k)
frame_vm_group_bin_16173 = frame (4k)
frame_vm_group_bin_16174 = frame (4k)
frame_vm_group_bin_16175 = frame (4k)
frame_vm_group_bin_16176 = frame (4k)
frame_vm_group_bin_16177 = frame (4k)
frame_vm_group_bin_16178 = frame (4k)
frame_vm_group_bin_16179 = frame (4k)
frame_vm_group_bin_1618 = frame (4k)
frame_vm_group_bin_16180 = frame (4k)
frame_vm_group_bin_16181 = frame (4k)
frame_vm_group_bin_16182 = frame (4k)
frame_vm_group_bin_16183 = frame (4k)
frame_vm_group_bin_16184 = frame (4k)
frame_vm_group_bin_16185 = frame (4k)
frame_vm_group_bin_16186 = frame (4k)
frame_vm_group_bin_16187 = frame (4k)
frame_vm_group_bin_16188 = frame (4k)
frame_vm_group_bin_16189 = frame (4k)
frame_vm_group_bin_1619 = frame (4k)
frame_vm_group_bin_16190 = frame (4k)
frame_vm_group_bin_16191 = frame (4k)
frame_vm_group_bin_16192 = frame (4k)
frame_vm_group_bin_16193 = frame (4k)
frame_vm_group_bin_16194 = frame (4k)
frame_vm_group_bin_16195 = frame (4k)
frame_vm_group_bin_16196 = frame (4k)
frame_vm_group_bin_16197 = frame (4k)
frame_vm_group_bin_16198 = frame (4k)
frame_vm_group_bin_16199 = frame (4k)
frame_vm_group_bin_1620 = frame (4k)
frame_vm_group_bin_16200 = frame (4k)
frame_vm_group_bin_16201 = frame (4k)
frame_vm_group_bin_16202 = frame (4k)
frame_vm_group_bin_16203 = frame (4k)
frame_vm_group_bin_16204 = frame (4k)
frame_vm_group_bin_16205 = frame (4k)
frame_vm_group_bin_16206 = frame (4k)
frame_vm_group_bin_16207 = frame (4k)
frame_vm_group_bin_16208 = frame (4k)
frame_vm_group_bin_16209 = frame (4k)
frame_vm_group_bin_1621 = frame (4k)
frame_vm_group_bin_16210 = frame (4k)
frame_vm_group_bin_16211 = frame (4k)
frame_vm_group_bin_16212 = frame (4k)
frame_vm_group_bin_16213 = frame (4k)
frame_vm_group_bin_16214 = frame (4k)
frame_vm_group_bin_16215 = frame (4k)
frame_vm_group_bin_16216 = frame (4k)
frame_vm_group_bin_16217 = frame (4k)
frame_vm_group_bin_16218 = frame (4k)
frame_vm_group_bin_16219 = frame (4k)
frame_vm_group_bin_1622 = frame (4k)
frame_vm_group_bin_16220 = frame (4k)
frame_vm_group_bin_16221 = frame (4k)
frame_vm_group_bin_16222 = frame (4k)
frame_vm_group_bin_16223 = frame (4k)
frame_vm_group_bin_16224 = frame (4k)
frame_vm_group_bin_16225 = frame (4k)
frame_vm_group_bin_16226 = frame (4k)
frame_vm_group_bin_16227 = frame (4k)
frame_vm_group_bin_16228 = frame (4k)
frame_vm_group_bin_16229 = frame (4k)
frame_vm_group_bin_1623 = frame (4k)
frame_vm_group_bin_16230 = frame (4k)
frame_vm_group_bin_16231 = frame (4k)
frame_vm_group_bin_16232 = frame (4k)
frame_vm_group_bin_16233 = frame (4k)
frame_vm_group_bin_16234 = frame (4k)
frame_vm_group_bin_16235 = frame (4k)
frame_vm_group_bin_16236 = frame (4k)
frame_vm_group_bin_16237 = frame (4k)
frame_vm_group_bin_16238 = frame (4k)
frame_vm_group_bin_16239 = frame (4k)
frame_vm_group_bin_1624 = frame (4k)
frame_vm_group_bin_16240 = frame (4k)
frame_vm_group_bin_16241 = frame (4k)
frame_vm_group_bin_16242 = frame (4k)
frame_vm_group_bin_16243 = frame (4k)
frame_vm_group_bin_16244 = frame (4k)
frame_vm_group_bin_16245 = frame (4k)
frame_vm_group_bin_16246 = frame (4k)
frame_vm_group_bin_16247 = frame (4k)
frame_vm_group_bin_16248 = frame (4k)
frame_vm_group_bin_16249 = frame (4k)
frame_vm_group_bin_1625 = frame (4k)
frame_vm_group_bin_16250 = frame (4k)
frame_vm_group_bin_16251 = frame (4k)
frame_vm_group_bin_16252 = frame (4k)
frame_vm_group_bin_16253 = frame (4k)
frame_vm_group_bin_16254 = frame (4k)
frame_vm_group_bin_16255 = frame (4k)
frame_vm_group_bin_16256 = frame (4k)
frame_vm_group_bin_16257 = frame (4k)
frame_vm_group_bin_16258 = frame (4k)
frame_vm_group_bin_16259 = frame (4k)
frame_vm_group_bin_1626 = frame (4k)
frame_vm_group_bin_16260 = frame (4k)
frame_vm_group_bin_16261 = frame (4k)
frame_vm_group_bin_16262 = frame (4k)
frame_vm_group_bin_16263 = frame (4k)
frame_vm_group_bin_16264 = frame (4k)
frame_vm_group_bin_16265 = frame (4k)
frame_vm_group_bin_16266 = frame (4k)
frame_vm_group_bin_16267 = frame (4k)
frame_vm_group_bin_16268 = frame (4k)
frame_vm_group_bin_16269 = frame (4k)
frame_vm_group_bin_1627 = frame (4k)
frame_vm_group_bin_16270 = frame (4k)
frame_vm_group_bin_16271 = frame (4k)
frame_vm_group_bin_16272 = frame (4k)
frame_vm_group_bin_16273 = frame (4k)
frame_vm_group_bin_16274 = frame (4k)
frame_vm_group_bin_16275 = frame (4k)
frame_vm_group_bin_16276 = frame (4k)
frame_vm_group_bin_16277 = frame (4k)
frame_vm_group_bin_16278 = frame (4k)
frame_vm_group_bin_16279 = frame (4k)
frame_vm_group_bin_1628 = frame (4k)
frame_vm_group_bin_16280 = frame (4k)
frame_vm_group_bin_16281 = frame (4k)
frame_vm_group_bin_16282 = frame (4k)
frame_vm_group_bin_16283 = frame (4k)
frame_vm_group_bin_16284 = frame (4k)
frame_vm_group_bin_16285 = frame (4k)
frame_vm_group_bin_16286 = frame (4k)
frame_vm_group_bin_16287 = frame (4k)
frame_vm_group_bin_16288 = frame (4k)
frame_vm_group_bin_16289 = frame (4k)
frame_vm_group_bin_1629 = frame (4k)
frame_vm_group_bin_16290 = frame (4k)
frame_vm_group_bin_16291 = frame (4k)
frame_vm_group_bin_16292 = frame (4k)
frame_vm_group_bin_16293 = frame (4k)
frame_vm_group_bin_16294 = frame (4k)
frame_vm_group_bin_16295 = frame (4k)
frame_vm_group_bin_16296 = frame (4k)
frame_vm_group_bin_16297 = frame (4k)
frame_vm_group_bin_16298 = frame (4k)
frame_vm_group_bin_16299 = frame (4k)
frame_vm_group_bin_1630 = frame (4k)
frame_vm_group_bin_16300 = frame (4k)
frame_vm_group_bin_16301 = frame (4k)
frame_vm_group_bin_16302 = frame (4k)
frame_vm_group_bin_16303 = frame (4k)
frame_vm_group_bin_16304 = frame (4k)
frame_vm_group_bin_16305 = frame (4k)
frame_vm_group_bin_16306 = frame (4k)
frame_vm_group_bin_16307 = frame (4k)
frame_vm_group_bin_16308 = frame (4k)
frame_vm_group_bin_16309 = frame (4k)
frame_vm_group_bin_1631 = frame (4k)
frame_vm_group_bin_16310 = frame (4k)
frame_vm_group_bin_16311 = frame (4k)
frame_vm_group_bin_16312 = frame (4k)
frame_vm_group_bin_16313 = frame (4k)
frame_vm_group_bin_16314 = frame (4k)
frame_vm_group_bin_16315 = frame (4k)
frame_vm_group_bin_16316 = frame (4k)
frame_vm_group_bin_16317 = frame (4k)
frame_vm_group_bin_16318 = frame (4k)
frame_vm_group_bin_16319 = frame (4k)
frame_vm_group_bin_1632 = frame (4k)
frame_vm_group_bin_16320 = frame (4k)
frame_vm_group_bin_16321 = frame (4k)
frame_vm_group_bin_16322 = frame (4k)
frame_vm_group_bin_16323 = frame (4k)
frame_vm_group_bin_16324 = frame (4k)
frame_vm_group_bin_16325 = frame (4k)
frame_vm_group_bin_16326 = frame (4k)
frame_vm_group_bin_16327 = frame (4k)
frame_vm_group_bin_16328 = frame (4k)
frame_vm_group_bin_16329 = frame (4k)
frame_vm_group_bin_16330 = frame (4k)
frame_vm_group_bin_16331 = frame (4k)
frame_vm_group_bin_16332 = frame (4k)
frame_vm_group_bin_16333 = frame (4k)
frame_vm_group_bin_16334 = frame (4k)
frame_vm_group_bin_16335 = frame (4k)
frame_vm_group_bin_16336 = frame (4k)
frame_vm_group_bin_16337 = frame (4k)
frame_vm_group_bin_16338 = frame (4k)
frame_vm_group_bin_16339 = frame (4k)
frame_vm_group_bin_1634 = frame (4k)
frame_vm_group_bin_16340 = frame (4k)
frame_vm_group_bin_16341 = frame (4k)
frame_vm_group_bin_16342 = frame (4k)
frame_vm_group_bin_16343 = frame (4k)
frame_vm_group_bin_16344 = frame (4k)
frame_vm_group_bin_16345 = frame (4k)
frame_vm_group_bin_16346 = frame (4k)
frame_vm_group_bin_16347 = frame (4k)
frame_vm_group_bin_16348 = frame (4k)
frame_vm_group_bin_16349 = frame (4k)
frame_vm_group_bin_1635 = frame (4k)
frame_vm_group_bin_16350 = frame (4k)
frame_vm_group_bin_16351 = frame (4k)
frame_vm_group_bin_16352 = frame (4k)
frame_vm_group_bin_16353 = frame (4k)
frame_vm_group_bin_16354 = frame (4k)
frame_vm_group_bin_16355 = frame (4k)
frame_vm_group_bin_16356 = frame (4k)
frame_vm_group_bin_16357 = frame (4k)
frame_vm_group_bin_16358 = frame (4k)
frame_vm_group_bin_16359 = frame (4k)
frame_vm_group_bin_1636 = frame (4k)
frame_vm_group_bin_16360 = frame (4k)
frame_vm_group_bin_16361 = frame (4k)
frame_vm_group_bin_16362 = frame (4k)
frame_vm_group_bin_16363 = frame (4k)
frame_vm_group_bin_16364 = frame (4k)
frame_vm_group_bin_16365 = frame (4k)
frame_vm_group_bin_16366 = frame (4k)
frame_vm_group_bin_16367 = frame (4k)
frame_vm_group_bin_16368 = frame (4k)
frame_vm_group_bin_16369 = frame (4k)
frame_vm_group_bin_1637 = frame (4k)
frame_vm_group_bin_16370 = frame (4k)
frame_vm_group_bin_16371 = frame (4k)
frame_vm_group_bin_16372 = frame (4k)
frame_vm_group_bin_16373 = frame (4k)
frame_vm_group_bin_16374 = frame (4k)
frame_vm_group_bin_16375 = frame (4k)
frame_vm_group_bin_16376 = frame (4k)
frame_vm_group_bin_16377 = frame (4k)
frame_vm_group_bin_16378 = frame (4k)
frame_vm_group_bin_16379 = frame (4k)
frame_vm_group_bin_1638 = frame (4k)
frame_vm_group_bin_16380 = frame (4k)
frame_vm_group_bin_16381 = frame (4k)
frame_vm_group_bin_16382 = frame (4k)
frame_vm_group_bin_16383 = frame (4k)
frame_vm_group_bin_16384 = frame (4k)
frame_vm_group_bin_16385 = frame (4k)
frame_vm_group_bin_16386 = frame (4k)
frame_vm_group_bin_16387 = frame (4k)
frame_vm_group_bin_16388 = frame (4k)
frame_vm_group_bin_16389 = frame (4k)
frame_vm_group_bin_1639 = frame (4k)
frame_vm_group_bin_16390 = frame (4k)
frame_vm_group_bin_16391 = frame (4k)
frame_vm_group_bin_16392 = frame (4k)
frame_vm_group_bin_16393 = frame (4k)
frame_vm_group_bin_16394 = frame (4k)
frame_vm_group_bin_16395 = frame (4k)
frame_vm_group_bin_16396 = frame (4k)
frame_vm_group_bin_16397 = frame (4k)
frame_vm_group_bin_16398 = frame (4k)
frame_vm_group_bin_16399 = frame (4k)
frame_vm_group_bin_1640 = frame (4k)
frame_vm_group_bin_16400 = frame (4k)
frame_vm_group_bin_16401 = frame (4k)
frame_vm_group_bin_16402 = frame (4k)
frame_vm_group_bin_16403 = frame (4k)
frame_vm_group_bin_16404 = frame (4k)
frame_vm_group_bin_16405 = frame (4k)
frame_vm_group_bin_16406 = frame (4k)
frame_vm_group_bin_16407 = frame (4k)
frame_vm_group_bin_16408 = frame (4k)
frame_vm_group_bin_16409 = frame (4k)
frame_vm_group_bin_1641 = frame (4k)
frame_vm_group_bin_16410 = frame (4k)
frame_vm_group_bin_16411 = frame (4k)
frame_vm_group_bin_16412 = frame (4k)
frame_vm_group_bin_16413 = frame (4k)
frame_vm_group_bin_16414 = frame (4k)
frame_vm_group_bin_16415 = frame (4k)
frame_vm_group_bin_16416 = frame (4k)
frame_vm_group_bin_16417 = frame (4k)
frame_vm_group_bin_16418 = frame (4k)
frame_vm_group_bin_16419 = frame (4k)
frame_vm_group_bin_1642 = frame (4k)
frame_vm_group_bin_16420 = frame (4k)
frame_vm_group_bin_16421 = frame (4k)
frame_vm_group_bin_16422 = frame (4k)
frame_vm_group_bin_16423 = frame (4k)
frame_vm_group_bin_16424 = frame (4k)
frame_vm_group_bin_16425 = frame (4k)
frame_vm_group_bin_16426 = frame (4k)
frame_vm_group_bin_16427 = frame (4k)
frame_vm_group_bin_16428 = frame (4k)
frame_vm_group_bin_16429 = frame (4k)
frame_vm_group_bin_1643 = frame (4k)
frame_vm_group_bin_16430 = frame (4k)
frame_vm_group_bin_16431 = frame (4k)
frame_vm_group_bin_16432 = frame (4k)
frame_vm_group_bin_16433 = frame (4k)
frame_vm_group_bin_16434 = frame (4k)
frame_vm_group_bin_16435 = frame (4k)
frame_vm_group_bin_16436 = frame (4k)
frame_vm_group_bin_16437 = frame (4k)
frame_vm_group_bin_16438 = frame (4k)
frame_vm_group_bin_16439 = frame (4k)
frame_vm_group_bin_1644 = frame (4k)
frame_vm_group_bin_16440 = frame (4k)
frame_vm_group_bin_16441 = frame (4k)
frame_vm_group_bin_16442 = frame (4k)
frame_vm_group_bin_16443 = frame (4k)
frame_vm_group_bin_16444 = frame (4k)
frame_vm_group_bin_16445 = frame (4k)
frame_vm_group_bin_16446 = frame (4k)
frame_vm_group_bin_16447 = frame (4k)
frame_vm_group_bin_16448 = frame (4k)
frame_vm_group_bin_16449 = frame (4k)
frame_vm_group_bin_1645 = frame (4k)
frame_vm_group_bin_16450 = frame (4k)
frame_vm_group_bin_16451 = frame (4k)
frame_vm_group_bin_16452 = frame (4k)
frame_vm_group_bin_16453 = frame (4k)
frame_vm_group_bin_16454 = frame (4k)
frame_vm_group_bin_16455 = frame (4k)
frame_vm_group_bin_16456 = frame (4k)
frame_vm_group_bin_16457 = frame (4k)
frame_vm_group_bin_16458 = frame (4k)
frame_vm_group_bin_16459 = frame (4k)
frame_vm_group_bin_1646 = frame (4k)
frame_vm_group_bin_16460 = frame (4k)
frame_vm_group_bin_16461 = frame (4k)
frame_vm_group_bin_16462 = frame (4k)
frame_vm_group_bin_16463 = frame (4k)
frame_vm_group_bin_16464 = frame (4k)
frame_vm_group_bin_16465 = frame (4k)
frame_vm_group_bin_16466 = frame (4k)
frame_vm_group_bin_16467 = frame (4k)
frame_vm_group_bin_16468 = frame (4k)
frame_vm_group_bin_16469 = frame (4k)
frame_vm_group_bin_1647 = frame (4k)
frame_vm_group_bin_16470 = frame (4k)
frame_vm_group_bin_16471 = frame (4k)
frame_vm_group_bin_16472 = frame (4k)
frame_vm_group_bin_16473 = frame (4k)
frame_vm_group_bin_16474 = frame (4k)
frame_vm_group_bin_16475 = frame (4k)
frame_vm_group_bin_16476 = frame (4k)
frame_vm_group_bin_16477 = frame (4k)
frame_vm_group_bin_16478 = frame (4k)
frame_vm_group_bin_16479 = frame (4k)
frame_vm_group_bin_1648 = frame (4k)
frame_vm_group_bin_16480 = frame (4k)
frame_vm_group_bin_16481 = frame (4k)
frame_vm_group_bin_16482 = frame (4k)
frame_vm_group_bin_16483 = frame (4k)
frame_vm_group_bin_16484 = frame (4k)
frame_vm_group_bin_16485 = frame (4k)
frame_vm_group_bin_16486 = frame (4k)
frame_vm_group_bin_16487 = frame (4k)
frame_vm_group_bin_16488 = frame (4k)
frame_vm_group_bin_16489 = frame (4k)
frame_vm_group_bin_1649 = frame (4k)
frame_vm_group_bin_16490 = frame (4k)
frame_vm_group_bin_16491 = frame (4k)
frame_vm_group_bin_16492 = frame (4k)
frame_vm_group_bin_16493 = frame (4k)
frame_vm_group_bin_16494 = frame (4k)
frame_vm_group_bin_16495 = frame (4k)
frame_vm_group_bin_16496 = frame (4k)
frame_vm_group_bin_16497 = frame (4k)
frame_vm_group_bin_16498 = frame (4k)
frame_vm_group_bin_16499 = frame (4k)
frame_vm_group_bin_1650 = frame (4k)
frame_vm_group_bin_16500 = frame (4k)
frame_vm_group_bin_16501 = frame (4k)
frame_vm_group_bin_16502 = frame (4k)
frame_vm_group_bin_16503 = frame (4k)
frame_vm_group_bin_16504 = frame (4k)
frame_vm_group_bin_16505 = frame (4k)
frame_vm_group_bin_16506 = frame (4k)
frame_vm_group_bin_16507 = frame (4k)
frame_vm_group_bin_16508 = frame (4k)
frame_vm_group_bin_16509 = frame (4k)
frame_vm_group_bin_1651 = frame (4k)
frame_vm_group_bin_16510 = frame (4k)
frame_vm_group_bin_16511 = frame (4k)
frame_vm_group_bin_16512 = frame (4k)
frame_vm_group_bin_16513 = frame (4k)
frame_vm_group_bin_16514 = frame (4k)
frame_vm_group_bin_16515 = frame (4k)
frame_vm_group_bin_16516 = frame (4k)
frame_vm_group_bin_16517 = frame (4k)
frame_vm_group_bin_16518 = frame (4k)
frame_vm_group_bin_16519 = frame (4k)
frame_vm_group_bin_1652 = frame (4k)
frame_vm_group_bin_16520 = frame (4k)
frame_vm_group_bin_16521 = frame (4k)
frame_vm_group_bin_16522 = frame (4k)
frame_vm_group_bin_16523 = frame (4k)
frame_vm_group_bin_16524 = frame (4k)
frame_vm_group_bin_16525 = frame (4k)
frame_vm_group_bin_16526 = frame (4k)
frame_vm_group_bin_16527 = frame (4k)
frame_vm_group_bin_16528 = frame (4k)
frame_vm_group_bin_16529 = frame (4k)
frame_vm_group_bin_1653 = frame (4k)
frame_vm_group_bin_16530 = frame (4k)
frame_vm_group_bin_16531 = frame (4k)
frame_vm_group_bin_16532 = frame (4k)
frame_vm_group_bin_16533 = frame (4k)
frame_vm_group_bin_16534 = frame (4k)
frame_vm_group_bin_16535 = frame (4k)
frame_vm_group_bin_16536 = frame (4k)
frame_vm_group_bin_16537 = frame (4k)
frame_vm_group_bin_16538 = frame (4k)
frame_vm_group_bin_16539 = frame (4k)
frame_vm_group_bin_1654 = frame (4k)
frame_vm_group_bin_16540 = frame (4k)
frame_vm_group_bin_16541 = frame (4k)
frame_vm_group_bin_16542 = frame (4k)
frame_vm_group_bin_16543 = frame (4k)
frame_vm_group_bin_16544 = frame (4k)
frame_vm_group_bin_16545 = frame (4k)
frame_vm_group_bin_16546 = frame (4k)
frame_vm_group_bin_16547 = frame (4k)
frame_vm_group_bin_16548 = frame (4k)
frame_vm_group_bin_16549 = frame (4k)
frame_vm_group_bin_1655 = frame (4k)
frame_vm_group_bin_16550 = frame (4k)
frame_vm_group_bin_16551 = frame (4k)
frame_vm_group_bin_16552 = frame (4k)
frame_vm_group_bin_16553 = frame (4k)
frame_vm_group_bin_16554 = frame (4k)
frame_vm_group_bin_16555 = frame (4k)
frame_vm_group_bin_16556 = frame (4k)
frame_vm_group_bin_16557 = frame (4k)
frame_vm_group_bin_16558 = frame (4k)
frame_vm_group_bin_16559 = frame (4k)
frame_vm_group_bin_1656 = frame (4k)
frame_vm_group_bin_16560 = frame (4k)
frame_vm_group_bin_16561 = frame (4k)
frame_vm_group_bin_16562 = frame (4k)
frame_vm_group_bin_16563 = frame (4k)
frame_vm_group_bin_16564 = frame (4k)
frame_vm_group_bin_16565 = frame (4k)
frame_vm_group_bin_16566 = frame (4k)
frame_vm_group_bin_16567 = frame (4k)
frame_vm_group_bin_16568 = frame (4k)
frame_vm_group_bin_16569 = frame (4k)
frame_vm_group_bin_1657 = frame (4k)
frame_vm_group_bin_16570 = frame (4k)
frame_vm_group_bin_16571 = frame (4k)
frame_vm_group_bin_16572 = frame (4k)
frame_vm_group_bin_16573 = frame (4k)
frame_vm_group_bin_16574 = frame (4k)
frame_vm_group_bin_16575 = frame (4k)
frame_vm_group_bin_16576 = frame (4k)
frame_vm_group_bin_16577 = frame (4k)
frame_vm_group_bin_16578 = frame (4k)
frame_vm_group_bin_16579 = frame (4k)
frame_vm_group_bin_1658 = frame (4k)
frame_vm_group_bin_16580 = frame (4k)
frame_vm_group_bin_16581 = frame (4k)
frame_vm_group_bin_16582 = frame (4k)
frame_vm_group_bin_16583 = frame (4k)
frame_vm_group_bin_16584 = frame (4k)
frame_vm_group_bin_16585 = frame (4k)
frame_vm_group_bin_16586 = frame (4k)
frame_vm_group_bin_16587 = frame (4k)
frame_vm_group_bin_16588 = frame (4k)
frame_vm_group_bin_16589 = frame (4k)
frame_vm_group_bin_1659 = frame (4k)
frame_vm_group_bin_16590 = frame (4k)
frame_vm_group_bin_16591 = frame (4k)
frame_vm_group_bin_16592 = frame (4k)
frame_vm_group_bin_16593 = frame (4k)
frame_vm_group_bin_16594 = frame (4k)
frame_vm_group_bin_16595 = frame (4k)
frame_vm_group_bin_16596 = frame (4k)
frame_vm_group_bin_16597 = frame (4k)
frame_vm_group_bin_16598 = frame (4k)
frame_vm_group_bin_16599 = frame (4k)
frame_vm_group_bin_1660 = frame (4k)
frame_vm_group_bin_16600 = frame (4k)
frame_vm_group_bin_16601 = frame (4k)
frame_vm_group_bin_16602 = frame (4k)
frame_vm_group_bin_16603 = frame (4k)
frame_vm_group_bin_16604 = frame (4k)
frame_vm_group_bin_16605 = frame (4k)
frame_vm_group_bin_16606 = frame (4k)
frame_vm_group_bin_16607 = frame (4k)
frame_vm_group_bin_16608 = frame (4k)
frame_vm_group_bin_16609 = frame (4k)
frame_vm_group_bin_1661 = frame (4k)
frame_vm_group_bin_16610 = frame (4k)
frame_vm_group_bin_16611 = frame (4k)
frame_vm_group_bin_16612 = frame (4k)
frame_vm_group_bin_16613 = frame (4k)
frame_vm_group_bin_16614 = frame (4k)
frame_vm_group_bin_16615 = frame (4k)
frame_vm_group_bin_16616 = frame (4k)
frame_vm_group_bin_16617 = frame (4k)
frame_vm_group_bin_16618 = frame (4k)
frame_vm_group_bin_16619 = frame (4k)
frame_vm_group_bin_1662 = frame (4k)
frame_vm_group_bin_16620 = frame (4k)
frame_vm_group_bin_16621 = frame (4k)
frame_vm_group_bin_16622 = frame (4k)
frame_vm_group_bin_16623 = frame (4k)
frame_vm_group_bin_16624 = frame (4k)
frame_vm_group_bin_16625 = frame (4k)
frame_vm_group_bin_16626 = frame (4k)
frame_vm_group_bin_16627 = frame (4k)
frame_vm_group_bin_16628 = frame (4k)
frame_vm_group_bin_16629 = frame (4k)
frame_vm_group_bin_1663 = frame (4k)
frame_vm_group_bin_16630 = frame (4k)
frame_vm_group_bin_16631 = frame (4k)
frame_vm_group_bin_16632 = frame (4k)
frame_vm_group_bin_16633 = frame (4k)
frame_vm_group_bin_16634 = frame (4k)
frame_vm_group_bin_16635 = frame (4k)
frame_vm_group_bin_16636 = frame (4k)
frame_vm_group_bin_16637 = frame (4k)
frame_vm_group_bin_16638 = frame (4k)
frame_vm_group_bin_16639 = frame (4k)
frame_vm_group_bin_1664 = frame (4k)
frame_vm_group_bin_16640 = frame (4k)
frame_vm_group_bin_16641 = frame (4k)
frame_vm_group_bin_16642 = frame (4k)
frame_vm_group_bin_16643 = frame (4k)
frame_vm_group_bin_16644 = frame (4k)
frame_vm_group_bin_16645 = frame (4k)
frame_vm_group_bin_16646 = frame (4k)
frame_vm_group_bin_16647 = frame (4k)
frame_vm_group_bin_16648 = frame (4k)
frame_vm_group_bin_16649 = frame (4k)
frame_vm_group_bin_1665 = frame (4k)
frame_vm_group_bin_16650 = frame (4k)
frame_vm_group_bin_16651 = frame (4k)
frame_vm_group_bin_16652 = frame (4k)
frame_vm_group_bin_16653 = frame (4k)
frame_vm_group_bin_16654 = frame (4k)
frame_vm_group_bin_16655 = frame (4k)
frame_vm_group_bin_16656 = frame (4k)
frame_vm_group_bin_16657 = frame (4k)
frame_vm_group_bin_16658 = frame (4k)
frame_vm_group_bin_16659 = frame (4k)
frame_vm_group_bin_16660 = frame (4k)
frame_vm_group_bin_16661 = frame (4k)
frame_vm_group_bin_16662 = frame (4k)
frame_vm_group_bin_16663 = frame (4k)
frame_vm_group_bin_16664 = frame (4k)
frame_vm_group_bin_16665 = frame (4k)
frame_vm_group_bin_16666 = frame (4k)
frame_vm_group_bin_16667 = frame (4k)
frame_vm_group_bin_16668 = frame (4k)
frame_vm_group_bin_16669 = frame (4k)
frame_vm_group_bin_1667 = frame (4k)
frame_vm_group_bin_16670 = frame (4k)
frame_vm_group_bin_16671 = frame (4k)
frame_vm_group_bin_16672 = frame (4k)
frame_vm_group_bin_16673 = frame (4k)
frame_vm_group_bin_16674 = frame (4k)
frame_vm_group_bin_16675 = frame (4k)
frame_vm_group_bin_16676 = frame (4k)
frame_vm_group_bin_16677 = frame (4k)
frame_vm_group_bin_16678 = frame (4k)
frame_vm_group_bin_16679 = frame (4k)
frame_vm_group_bin_1668 = frame (4k)
frame_vm_group_bin_16680 = frame (4k)
frame_vm_group_bin_16681 = frame (4k)
frame_vm_group_bin_16682 = frame (4k)
frame_vm_group_bin_16683 = frame (4k)
frame_vm_group_bin_16684 = frame (4k)
frame_vm_group_bin_16685 = frame (4k)
frame_vm_group_bin_16686 = frame (4k)
frame_vm_group_bin_16687 = frame (4k)
frame_vm_group_bin_16688 = frame (4k)
frame_vm_group_bin_16689 = frame (4k)
frame_vm_group_bin_1669 = frame (4k)
frame_vm_group_bin_16690 = frame (4k)
frame_vm_group_bin_16691 = frame (4k)
frame_vm_group_bin_16692 = frame (4k)
frame_vm_group_bin_16693 = frame (4k)
frame_vm_group_bin_16694 = frame (4k)
frame_vm_group_bin_16695 = frame (4k)
frame_vm_group_bin_16696 = frame (4k)
frame_vm_group_bin_16697 = frame (4k)
frame_vm_group_bin_16698 = frame (4k)
frame_vm_group_bin_16699 = frame (4k)
frame_vm_group_bin_1670 = frame (4k)
frame_vm_group_bin_16700 = frame (4k)
frame_vm_group_bin_16701 = frame (4k)
frame_vm_group_bin_16702 = frame (4k)
frame_vm_group_bin_16703 = frame (4k)
frame_vm_group_bin_16704 = frame (4k)
frame_vm_group_bin_16705 = frame (4k)
frame_vm_group_bin_16706 = frame (4k)
frame_vm_group_bin_16707 = frame (4k)
frame_vm_group_bin_16708 = frame (4k)
frame_vm_group_bin_16709 = frame (4k)
frame_vm_group_bin_1671 = frame (4k)
frame_vm_group_bin_16710 = frame (4k)
frame_vm_group_bin_16711 = frame (4k)
frame_vm_group_bin_16712 = frame (4k)
frame_vm_group_bin_16713 = frame (4k)
frame_vm_group_bin_16714 = frame (4k)
frame_vm_group_bin_16715 = frame (4k)
frame_vm_group_bin_16716 = frame (4k)
frame_vm_group_bin_16717 = frame (4k)
frame_vm_group_bin_16718 = frame (4k)
frame_vm_group_bin_16719 = frame (4k)
frame_vm_group_bin_1672 = frame (4k)
frame_vm_group_bin_16720 = frame (4k)
frame_vm_group_bin_16721 = frame (4k)
frame_vm_group_bin_16722 = frame (4k)
frame_vm_group_bin_16723 = frame (4k)
frame_vm_group_bin_16724 = frame (4k)
frame_vm_group_bin_16725 = frame (4k)
frame_vm_group_bin_16726 = frame (4k)
frame_vm_group_bin_16727 = frame (4k)
frame_vm_group_bin_16728 = frame (4k)
frame_vm_group_bin_16729 = frame (4k)
frame_vm_group_bin_1673 = frame (4k)
frame_vm_group_bin_16730 = frame (4k)
frame_vm_group_bin_16731 = frame (4k)
frame_vm_group_bin_16732 = frame (4k)
frame_vm_group_bin_16733 = frame (4k)
frame_vm_group_bin_16734 = frame (4k)
frame_vm_group_bin_16735 = frame (4k)
frame_vm_group_bin_16736 = frame (4k)
frame_vm_group_bin_16737 = frame (4k)
frame_vm_group_bin_16738 = frame (4k)
frame_vm_group_bin_16739 = frame (4k)
frame_vm_group_bin_1674 = frame (4k)
frame_vm_group_bin_16740 = frame (4k)
frame_vm_group_bin_16741 = frame (4k)
frame_vm_group_bin_16742 = frame (4k)
frame_vm_group_bin_16743 = frame (4k)
frame_vm_group_bin_16744 = frame (4k)
frame_vm_group_bin_16745 = frame (4k)
frame_vm_group_bin_16746 = frame (4k)
frame_vm_group_bin_16747 = frame (4k)
frame_vm_group_bin_16748 = frame (4k)
frame_vm_group_bin_16749 = frame (4k)
frame_vm_group_bin_1675 = frame (4k)
frame_vm_group_bin_16750 = frame (4k)
frame_vm_group_bin_16751 = frame (4k)
frame_vm_group_bin_16752 = frame (4k)
frame_vm_group_bin_16753 = frame (4k)
frame_vm_group_bin_16754 = frame (4k)
frame_vm_group_bin_16755 = frame (4k)
frame_vm_group_bin_16756 = frame (4k)
frame_vm_group_bin_16757 = frame (4k)
frame_vm_group_bin_16758 = frame (4k)
frame_vm_group_bin_16759 = frame (4k)
frame_vm_group_bin_1676 = frame (4k)
frame_vm_group_bin_16760 = frame (4k)
frame_vm_group_bin_16761 = frame (4k)
frame_vm_group_bin_16762 = frame (4k)
frame_vm_group_bin_16763 = frame (4k)
frame_vm_group_bin_16764 = frame (4k)
frame_vm_group_bin_16765 = frame (4k)
frame_vm_group_bin_16766 = frame (4k)
frame_vm_group_bin_16767 = frame (4k)
frame_vm_group_bin_16768 = frame (4k)
frame_vm_group_bin_16769 = frame (4k)
frame_vm_group_bin_1677 = frame (4k)
frame_vm_group_bin_16770 = frame (4k)
frame_vm_group_bin_16771 = frame (4k)
frame_vm_group_bin_16772 = frame (4k)
frame_vm_group_bin_16773 = frame (4k)
frame_vm_group_bin_16774 = frame (4k)
frame_vm_group_bin_16775 = frame (4k)
frame_vm_group_bin_16776 = frame (4k)
frame_vm_group_bin_16777 = frame (4k)
frame_vm_group_bin_16778 = frame (4k)
frame_vm_group_bin_16779 = frame (4k)
frame_vm_group_bin_1678 = frame (4k)
frame_vm_group_bin_16780 = frame (4k)
frame_vm_group_bin_16781 = frame (4k)
frame_vm_group_bin_16782 = frame (4k)
frame_vm_group_bin_16783 = frame (4k)
frame_vm_group_bin_16784 = frame (4k)
frame_vm_group_bin_16785 = frame (4k)
frame_vm_group_bin_16786 = frame (4k)
frame_vm_group_bin_16787 = frame (4k)
frame_vm_group_bin_16788 = frame (4k)
frame_vm_group_bin_16789 = frame (4k)
frame_vm_group_bin_1679 = frame (4k)
frame_vm_group_bin_16790 = frame (4k)
frame_vm_group_bin_16791 = frame (4k)
frame_vm_group_bin_16792 = frame (4k)
frame_vm_group_bin_16793 = frame (4k)
frame_vm_group_bin_16794 = frame (4k)
frame_vm_group_bin_16795 = frame (4k)
frame_vm_group_bin_16796 = frame (4k)
frame_vm_group_bin_16797 = frame (4k)
frame_vm_group_bin_16798 = frame (4k)
frame_vm_group_bin_16799 = frame (4k)
frame_vm_group_bin_1680 = frame (4k)
frame_vm_group_bin_16800 = frame (4k)
frame_vm_group_bin_16801 = frame (4k)
frame_vm_group_bin_16802 = frame (4k)
frame_vm_group_bin_16803 = frame (4k)
frame_vm_group_bin_16804 = frame (4k)
frame_vm_group_bin_16805 = frame (4k)
frame_vm_group_bin_16806 = frame (4k)
frame_vm_group_bin_16807 = frame (4k)
frame_vm_group_bin_16808 = frame (4k)
frame_vm_group_bin_16809 = frame (4k)
frame_vm_group_bin_1681 = frame (4k)
frame_vm_group_bin_16810 = frame (4k)
frame_vm_group_bin_16811 = frame (4k)
frame_vm_group_bin_16812 = frame (4k)
frame_vm_group_bin_16813 = frame (4k)
frame_vm_group_bin_16814 = frame (4k)
frame_vm_group_bin_16815 = frame (4k)
frame_vm_group_bin_16816 = frame (4k)
frame_vm_group_bin_16817 = frame (4k)
frame_vm_group_bin_16818 = frame (4k)
frame_vm_group_bin_16819 = frame (4k)
frame_vm_group_bin_1682 = frame (4k)
frame_vm_group_bin_16820 = frame (4k)
frame_vm_group_bin_16821 = frame (4k)
frame_vm_group_bin_16822 = frame (4k)
frame_vm_group_bin_16823 = frame (4k)
frame_vm_group_bin_16824 = frame (4k)
frame_vm_group_bin_16825 = frame (4k)
frame_vm_group_bin_16826 = frame (4k)
frame_vm_group_bin_16827 = frame (4k)
frame_vm_group_bin_16828 = frame (4k)
frame_vm_group_bin_16829 = frame (4k)
frame_vm_group_bin_1683 = frame (4k)
frame_vm_group_bin_16830 = frame (4k)
frame_vm_group_bin_16831 = frame (4k)
frame_vm_group_bin_16832 = frame (4k)
frame_vm_group_bin_16833 = frame (4k)
frame_vm_group_bin_16834 = frame (4k)
frame_vm_group_bin_16835 = frame (4k)
frame_vm_group_bin_16836 = frame (4k)
frame_vm_group_bin_16837 = frame (4k)
frame_vm_group_bin_16838 = frame (4k)
frame_vm_group_bin_16839 = frame (4k)
frame_vm_group_bin_1684 = frame (4k)
frame_vm_group_bin_16840 = frame (4k)
frame_vm_group_bin_16841 = frame (4k)
frame_vm_group_bin_16842 = frame (4k)
frame_vm_group_bin_16843 = frame (4k)
frame_vm_group_bin_16844 = frame (4k)
frame_vm_group_bin_16845 = frame (4k)
frame_vm_group_bin_16846 = frame (4k)
frame_vm_group_bin_16847 = frame (4k)
frame_vm_group_bin_16848 = frame (4k)
frame_vm_group_bin_16849 = frame (4k)
frame_vm_group_bin_1685 = frame (4k)
frame_vm_group_bin_16850 = frame (4k)
frame_vm_group_bin_16851 = frame (4k)
frame_vm_group_bin_16852 = frame (4k)
frame_vm_group_bin_16853 = frame (4k)
frame_vm_group_bin_16854 = frame (4k)
frame_vm_group_bin_16855 = frame (4k)
frame_vm_group_bin_16856 = frame (4k)
frame_vm_group_bin_16857 = frame (4k)
frame_vm_group_bin_16858 = frame (4k)
frame_vm_group_bin_16859 = frame (4k)
frame_vm_group_bin_1686 = frame (4k)
frame_vm_group_bin_16860 = frame (4k)
frame_vm_group_bin_16861 = frame (4k)
frame_vm_group_bin_16862 = frame (4k)
frame_vm_group_bin_16863 = frame (4k)
frame_vm_group_bin_16864 = frame (4k)
frame_vm_group_bin_16865 = frame (4k)
frame_vm_group_bin_16866 = frame (4k)
frame_vm_group_bin_16867 = frame (4k)
frame_vm_group_bin_16868 = frame (4k)
frame_vm_group_bin_16869 = frame (4k)
frame_vm_group_bin_1687 = frame (4k)
frame_vm_group_bin_16870 = frame (4k)
frame_vm_group_bin_16871 = frame (4k)
frame_vm_group_bin_16872 = frame (4k)
frame_vm_group_bin_16873 = frame (4k)
frame_vm_group_bin_16874 = frame (4k)
frame_vm_group_bin_16875 = frame (4k)
frame_vm_group_bin_16876 = frame (4k)
frame_vm_group_bin_16877 = frame (4k)
frame_vm_group_bin_16878 = frame (4k)
frame_vm_group_bin_16879 = frame (4k)
frame_vm_group_bin_1688 = frame (4k)
frame_vm_group_bin_16880 = frame (4k)
frame_vm_group_bin_16881 = frame (4k)
frame_vm_group_bin_16882 = frame (4k)
frame_vm_group_bin_16883 = frame (4k)
frame_vm_group_bin_16884 = frame (4k)
frame_vm_group_bin_16885 = frame (4k)
frame_vm_group_bin_16886 = frame (4k)
frame_vm_group_bin_16887 = frame (4k)
frame_vm_group_bin_16888 = frame (4k)
frame_vm_group_bin_16889 = frame (4k)
frame_vm_group_bin_1689 = frame (4k)
frame_vm_group_bin_16890 = frame (4k)
frame_vm_group_bin_16891 = frame (4k)
frame_vm_group_bin_16892 = frame (4k)
frame_vm_group_bin_16893 = frame (4k)
frame_vm_group_bin_16894 = frame (4k)
frame_vm_group_bin_16895 = frame (4k)
frame_vm_group_bin_16896 = frame (4k)
frame_vm_group_bin_16897 = frame (4k)
frame_vm_group_bin_16898 = frame (4k)
frame_vm_group_bin_16899 = frame (4k)
frame_vm_group_bin_1690 = frame (4k)
frame_vm_group_bin_16900 = frame (4k)
frame_vm_group_bin_16901 = frame (4k)
frame_vm_group_bin_16902 = frame (4k)
frame_vm_group_bin_16903 = frame (4k)
frame_vm_group_bin_16904 = frame (4k)
frame_vm_group_bin_16905 = frame (4k)
frame_vm_group_bin_16906 = frame (4k)
frame_vm_group_bin_16907 = frame (4k)
frame_vm_group_bin_16908 = frame (4k)
frame_vm_group_bin_16909 = frame (4k)
frame_vm_group_bin_1691 = frame (4k)
frame_vm_group_bin_16910 = frame (4k)
frame_vm_group_bin_16911 = frame (4k)
frame_vm_group_bin_16912 = frame (4k)
frame_vm_group_bin_16913 = frame (4k)
frame_vm_group_bin_16914 = frame (4k)
frame_vm_group_bin_16915 = frame (4k)
frame_vm_group_bin_16916 = frame (4k)
frame_vm_group_bin_16917 = frame (4k)
frame_vm_group_bin_16918 = frame (4k)
frame_vm_group_bin_16919 = frame (4k)
frame_vm_group_bin_1692 = frame (4k)
frame_vm_group_bin_16920 = frame (4k)
frame_vm_group_bin_16921 = frame (4k)
frame_vm_group_bin_16922 = frame (4k)
frame_vm_group_bin_16923 = frame (4k)
frame_vm_group_bin_16924 = frame (4k)
frame_vm_group_bin_16925 = frame (4k)
frame_vm_group_bin_16926 = frame (4k)
frame_vm_group_bin_16927 = frame (4k)
frame_vm_group_bin_16928 = frame (4k)
frame_vm_group_bin_16929 = frame (4k)
frame_vm_group_bin_1693 = frame (4k)
frame_vm_group_bin_16930 = frame (4k)
frame_vm_group_bin_16931 = frame (4k)
frame_vm_group_bin_16932 = frame (4k)
frame_vm_group_bin_16933 = frame (4k)
frame_vm_group_bin_16934 = frame (4k)
frame_vm_group_bin_16935 = frame (4k)
frame_vm_group_bin_16936 = frame (4k)
frame_vm_group_bin_16937 = frame (4k)
frame_vm_group_bin_16938 = frame (4k)
frame_vm_group_bin_16939 = frame (4k)
frame_vm_group_bin_1694 = frame (4k)
frame_vm_group_bin_16940 = frame (4k)
frame_vm_group_bin_16941 = frame (4k)
frame_vm_group_bin_16942 = frame (4k)
frame_vm_group_bin_16943 = frame (4k)
frame_vm_group_bin_16944 = frame (4k)
frame_vm_group_bin_16945 = frame (4k)
frame_vm_group_bin_16946 = frame (4k)
frame_vm_group_bin_16947 = frame (4k)
frame_vm_group_bin_16948 = frame (4k)
frame_vm_group_bin_16949 = frame (4k)
frame_vm_group_bin_1695 = frame (4k)
frame_vm_group_bin_16950 = frame (4k)
frame_vm_group_bin_16951 = frame (4k)
frame_vm_group_bin_16952 = frame (4k)
frame_vm_group_bin_16953 = frame (4k)
frame_vm_group_bin_16954 = frame (4k)
frame_vm_group_bin_16955 = frame (4k)
frame_vm_group_bin_16956 = frame (4k)
frame_vm_group_bin_16957 = frame (4k)
frame_vm_group_bin_16958 = frame (4k)
frame_vm_group_bin_16959 = frame (4k)
frame_vm_group_bin_1696 = frame (4k)
frame_vm_group_bin_16960 = frame (4k)
frame_vm_group_bin_16961 = frame (4k)
frame_vm_group_bin_16962 = frame (4k)
frame_vm_group_bin_16963 = frame (4k)
frame_vm_group_bin_16964 = frame (4k)
frame_vm_group_bin_16965 = frame (4k)
frame_vm_group_bin_16966 = frame (4k)
frame_vm_group_bin_16967 = frame (4k)
frame_vm_group_bin_16968 = frame (4k)
frame_vm_group_bin_16969 = frame (4k)
frame_vm_group_bin_1697 = frame (4k)
frame_vm_group_bin_16970 = frame (4k)
frame_vm_group_bin_16971 = frame (4k)
frame_vm_group_bin_16972 = frame (4k)
frame_vm_group_bin_16973 = frame (4k)
frame_vm_group_bin_16974 = frame (4k)
frame_vm_group_bin_16975 = frame (4k)
frame_vm_group_bin_16976 = frame (4k)
frame_vm_group_bin_16977 = frame (4k)
frame_vm_group_bin_16978 = frame (4k)
frame_vm_group_bin_16979 = frame (4k)
frame_vm_group_bin_1698 = frame (4k)
frame_vm_group_bin_16980 = frame (4k)
frame_vm_group_bin_16981 = frame (4k)
frame_vm_group_bin_16982 = frame (4k)
frame_vm_group_bin_16983 = frame (4k)
frame_vm_group_bin_16984 = frame (4k)
frame_vm_group_bin_16985 = frame (4k)
frame_vm_group_bin_16986 = frame (4k)
frame_vm_group_bin_16987 = frame (4k)
frame_vm_group_bin_16988 = frame (4k)
frame_vm_group_bin_16989 = frame (4k)
frame_vm_group_bin_1699 = frame (4k)
frame_vm_group_bin_16990 = frame (4k)
frame_vm_group_bin_16991 = frame (4k)
frame_vm_group_bin_16992 = frame (4k)
frame_vm_group_bin_16993 = frame (4k)
frame_vm_group_bin_16994 = frame (4k)
frame_vm_group_bin_16995 = frame (4k)
frame_vm_group_bin_16996 = frame (4k)
frame_vm_group_bin_16997 = frame (4k)
frame_vm_group_bin_16998 = frame (4k)
frame_vm_group_bin_16999 = frame (4k)
frame_vm_group_bin_1700 = frame (4k)
frame_vm_group_bin_17000 = frame (4k)
frame_vm_group_bin_17001 = frame (4k)
frame_vm_group_bin_17002 = frame (4k)
frame_vm_group_bin_17003 = frame (4k)
frame_vm_group_bin_17004 = frame (4k)
frame_vm_group_bin_17005 = frame (4k)
frame_vm_group_bin_17006 = frame (4k)
frame_vm_group_bin_17007 = frame (4k)
frame_vm_group_bin_17008 = frame (4k)
frame_vm_group_bin_17009 = frame (4k)
frame_vm_group_bin_1701 = frame (4k)
frame_vm_group_bin_17010 = frame (4k)
frame_vm_group_bin_17011 = frame (4k)
frame_vm_group_bin_17012 = frame (4k)
frame_vm_group_bin_17013 = frame (4k)
frame_vm_group_bin_17014 = frame (4k)
frame_vm_group_bin_17015 = frame (4k)
frame_vm_group_bin_17016 = frame (4k)
frame_vm_group_bin_17017 = frame (4k)
frame_vm_group_bin_17018 = frame (4k)
frame_vm_group_bin_17019 = frame (4k)
frame_vm_group_bin_1702 = frame (4k)
frame_vm_group_bin_17020 = frame (4k)
frame_vm_group_bin_17021 = frame (4k)
frame_vm_group_bin_17022 = frame (4k)
frame_vm_group_bin_17023 = frame (4k)
frame_vm_group_bin_17024 = frame (4k)
frame_vm_group_bin_17025 = frame (4k)
frame_vm_group_bin_17026 = frame (4k)
frame_vm_group_bin_17027 = frame (4k)
frame_vm_group_bin_17028 = frame (4k)
frame_vm_group_bin_17029 = frame (4k)
frame_vm_group_bin_1703 = frame (4k)
frame_vm_group_bin_17030 = frame (4k)
frame_vm_group_bin_17031 = frame (4k)
frame_vm_group_bin_17032 = frame (4k)
frame_vm_group_bin_17033 = frame (4k)
frame_vm_group_bin_17034 = frame (4k)
frame_vm_group_bin_17035 = frame (4k)
frame_vm_group_bin_17036 = frame (4k)
frame_vm_group_bin_17037 = frame (4k)
frame_vm_group_bin_17038 = frame (4k)
frame_vm_group_bin_17039 = frame (4k)
frame_vm_group_bin_1704 = frame (4k)
frame_vm_group_bin_17040 = frame (4k)
frame_vm_group_bin_17041 = frame (4k)
frame_vm_group_bin_17042 = frame (4k)
frame_vm_group_bin_17043 = frame (4k)
frame_vm_group_bin_17044 = frame (4k)
frame_vm_group_bin_17045 = frame (4k)
frame_vm_group_bin_17046 = frame (4k)
frame_vm_group_bin_17047 = frame (4k)
frame_vm_group_bin_17048 = frame (4k)
frame_vm_group_bin_17049 = frame (4k)
frame_vm_group_bin_1705 = frame (4k)
frame_vm_group_bin_17050 = frame (4k)
frame_vm_group_bin_17051 = frame (4k)
frame_vm_group_bin_17052 = frame (4k)
frame_vm_group_bin_17053 = frame (4k)
frame_vm_group_bin_17054 = frame (4k)
frame_vm_group_bin_17055 = frame (4k)
frame_vm_group_bin_17056 = frame (4k)
frame_vm_group_bin_17057 = frame (4k)
frame_vm_group_bin_17058 = frame (4k)
frame_vm_group_bin_17059 = frame (4k)
frame_vm_group_bin_1706 = frame (4k)
frame_vm_group_bin_17060 = frame (4k)
frame_vm_group_bin_17061 = frame (4k)
frame_vm_group_bin_17062 = frame (4k)
frame_vm_group_bin_17063 = frame (4k)
frame_vm_group_bin_17064 = frame (4k)
frame_vm_group_bin_17065 = frame (4k)
frame_vm_group_bin_17066 = frame (4k)
frame_vm_group_bin_17067 = frame (4k)
frame_vm_group_bin_17068 = frame (4k)
frame_vm_group_bin_17069 = frame (4k)
frame_vm_group_bin_1707 = frame (4k)
frame_vm_group_bin_17070 = frame (4k)
frame_vm_group_bin_17071 = frame (4k)
frame_vm_group_bin_17072 = frame (4k)
frame_vm_group_bin_17073 = frame (4k)
frame_vm_group_bin_17074 = frame (4k)
frame_vm_group_bin_17075 = frame (4k)
frame_vm_group_bin_17076 = frame (4k)
frame_vm_group_bin_17077 = frame (4k)
frame_vm_group_bin_17078 = frame (4k)
frame_vm_group_bin_17079 = frame (4k)
frame_vm_group_bin_1708 = frame (4k)
frame_vm_group_bin_17080 = frame (4k)
frame_vm_group_bin_17081 = frame (4k)
frame_vm_group_bin_17082 = frame (4k)
frame_vm_group_bin_17083 = frame (4k)
frame_vm_group_bin_17084 = frame (4k)
frame_vm_group_bin_17085 = frame (4k)
frame_vm_group_bin_17086 = frame (4k)
frame_vm_group_bin_17087 = frame (4k)
frame_vm_group_bin_17088 = frame (4k)
frame_vm_group_bin_17089 = frame (4k)
frame_vm_group_bin_1709 = frame (4k)
frame_vm_group_bin_17090 = frame (4k)
frame_vm_group_bin_17091 = frame (4k)
frame_vm_group_bin_17092 = frame (4k)
frame_vm_group_bin_17093 = frame (4k)
frame_vm_group_bin_17094 = frame (4k)
frame_vm_group_bin_17095 = frame (4k)
frame_vm_group_bin_17096 = frame (4k)
frame_vm_group_bin_17097 = frame (4k)
frame_vm_group_bin_17098 = frame (4k)
frame_vm_group_bin_17099 = frame (4k)
frame_vm_group_bin_1710 = frame (4k)
frame_vm_group_bin_17100 = frame (4k)
frame_vm_group_bin_17101 = frame (4k)
frame_vm_group_bin_17102 = frame (4k)
frame_vm_group_bin_17103 = frame (4k)
frame_vm_group_bin_17104 = frame (4k)
frame_vm_group_bin_17105 = frame (4k)
frame_vm_group_bin_17106 = frame (4k)
frame_vm_group_bin_17107 = frame (4k)
frame_vm_group_bin_17108 = frame (4k)
frame_vm_group_bin_17109 = frame (4k)
frame_vm_group_bin_1711 = frame (4k)
frame_vm_group_bin_17110 = frame (4k)
frame_vm_group_bin_17111 = frame (4k)
frame_vm_group_bin_17112 = frame (4k)
frame_vm_group_bin_17113 = frame (4k)
frame_vm_group_bin_17114 = frame (4k)
frame_vm_group_bin_17115 = frame (4k)
frame_vm_group_bin_17116 = frame (4k)
frame_vm_group_bin_17117 = frame (4k)
frame_vm_group_bin_17118 = frame (4k)
frame_vm_group_bin_17119 = frame (4k)
frame_vm_group_bin_1712 = frame (4k)
frame_vm_group_bin_17120 = frame (4k)
frame_vm_group_bin_17121 = frame (4k)
frame_vm_group_bin_17122 = frame (4k)
frame_vm_group_bin_17123 = frame (4k)
frame_vm_group_bin_17124 = frame (4k)
frame_vm_group_bin_17125 = frame (4k)
frame_vm_group_bin_17126 = frame (4k)
frame_vm_group_bin_17127 = frame (4k)
frame_vm_group_bin_17128 = frame (4k)
frame_vm_group_bin_17129 = frame (4k)
frame_vm_group_bin_1713 = frame (4k)
frame_vm_group_bin_17130 = frame (4k)
frame_vm_group_bin_17131 = frame (4k)
frame_vm_group_bin_17132 = frame (4k)
frame_vm_group_bin_17133 = frame (4k)
frame_vm_group_bin_17134 = frame (4k)
frame_vm_group_bin_17135 = frame (4k)
frame_vm_group_bin_17136 = frame (4k)
frame_vm_group_bin_17137 = frame (4k)
frame_vm_group_bin_17138 = frame (4k)
frame_vm_group_bin_17139 = frame (4k)
frame_vm_group_bin_1714 = frame (4k)
frame_vm_group_bin_17140 = frame (4k)
frame_vm_group_bin_17141 = frame (4k)
frame_vm_group_bin_17142 = frame (4k)
frame_vm_group_bin_17143 = frame (4k)
frame_vm_group_bin_17144 = frame (4k)
frame_vm_group_bin_17145 = frame (4k)
frame_vm_group_bin_17146 = frame (4k)
frame_vm_group_bin_17147 = frame (4k)
frame_vm_group_bin_17148 = frame (4k)
frame_vm_group_bin_17149 = frame (4k)
frame_vm_group_bin_1715 = frame (4k)
frame_vm_group_bin_17150 = frame (4k)
frame_vm_group_bin_17151 = frame (4k)
frame_vm_group_bin_17152 = frame (4k)
frame_vm_group_bin_17153 = frame (4k)
frame_vm_group_bin_17154 = frame (4k)
frame_vm_group_bin_17155 = frame (4k)
frame_vm_group_bin_17156 = frame (4k)
frame_vm_group_bin_17157 = frame (4k)
frame_vm_group_bin_17158 = frame (4k)
frame_vm_group_bin_17159 = frame (4k)
frame_vm_group_bin_1716 = frame (4k)
frame_vm_group_bin_17160 = frame (4k)
frame_vm_group_bin_17161 = frame (4k)
frame_vm_group_bin_17162 = frame (4k)
frame_vm_group_bin_17163 = frame (4k)
frame_vm_group_bin_17164 = frame (4k)
frame_vm_group_bin_17165 = frame (4k)
frame_vm_group_bin_17166 = frame (4k)
frame_vm_group_bin_17167 = frame (4k)
frame_vm_group_bin_17168 = frame (4k)
frame_vm_group_bin_17169 = frame (4k)
frame_vm_group_bin_1717 = frame (4k)
frame_vm_group_bin_17170 = frame (4k)
frame_vm_group_bin_17171 = frame (4k)
frame_vm_group_bin_17172 = frame (4k)
frame_vm_group_bin_17173 = frame (4k)
frame_vm_group_bin_17174 = frame (4k)
frame_vm_group_bin_17175 = frame (4k)
frame_vm_group_bin_17176 = frame (4k)
frame_vm_group_bin_17177 = frame (4k)
frame_vm_group_bin_17178 = frame (4k)
frame_vm_group_bin_17179 = frame (4k)
frame_vm_group_bin_1718 = frame (4k)
frame_vm_group_bin_17180 = frame (4k)
frame_vm_group_bin_17181 = frame (4k)
frame_vm_group_bin_17182 = frame (4k)
frame_vm_group_bin_17183 = frame (4k)
frame_vm_group_bin_17184 = frame (4k)
frame_vm_group_bin_17185 = frame (4k)
frame_vm_group_bin_17186 = frame (4k)
frame_vm_group_bin_17187 = frame (4k)
frame_vm_group_bin_17188 = frame (4k)
frame_vm_group_bin_17189 = frame (4k)
frame_vm_group_bin_1719 = frame (4k)
frame_vm_group_bin_17190 = frame (4k)
frame_vm_group_bin_17191 = frame (4k)
frame_vm_group_bin_17192 = frame (4k)
frame_vm_group_bin_17193 = frame (4k)
frame_vm_group_bin_17194 = frame (4k)
frame_vm_group_bin_17195 = frame (4k)
frame_vm_group_bin_17196 = frame (4k)
frame_vm_group_bin_17197 = frame (4k)
frame_vm_group_bin_17198 = frame (4k)
frame_vm_group_bin_17199 = frame (4k)
frame_vm_group_bin_1720 = frame (4k)
frame_vm_group_bin_17200 = frame (4k)
frame_vm_group_bin_17201 = frame (4k)
frame_vm_group_bin_17202 = frame (4k)
frame_vm_group_bin_17203 = frame (4k)
frame_vm_group_bin_17204 = frame (4k)
frame_vm_group_bin_17205 = frame (4k)
frame_vm_group_bin_17206 = frame (4k)
frame_vm_group_bin_17207 = frame (4k)
frame_vm_group_bin_17208 = frame (4k)
frame_vm_group_bin_17209 = frame (4k)
frame_vm_group_bin_1721 = frame (4k)
frame_vm_group_bin_17210 = frame (4k)
frame_vm_group_bin_17211 = frame (4k)
frame_vm_group_bin_17212 = frame (4k)
frame_vm_group_bin_17213 = frame (4k)
frame_vm_group_bin_17214 = frame (4k)
frame_vm_group_bin_17215 = frame (4k)
frame_vm_group_bin_17216 = frame (4k)
frame_vm_group_bin_17217 = frame (4k)
frame_vm_group_bin_17218 = frame (4k)
frame_vm_group_bin_17219 = frame (4k)
frame_vm_group_bin_1722 = frame (4k)
frame_vm_group_bin_17220 = frame (4k)
frame_vm_group_bin_17221 = frame (4k)
frame_vm_group_bin_17222 = frame (4k)
frame_vm_group_bin_17223 = frame (4k)
frame_vm_group_bin_17224 = frame (4k)
frame_vm_group_bin_17225 = frame (4k)
frame_vm_group_bin_17226 = frame (4k)
frame_vm_group_bin_17227 = frame (4k)
frame_vm_group_bin_17228 = frame (4k)
frame_vm_group_bin_17229 = frame (4k)
frame_vm_group_bin_1723 = frame (4k)
frame_vm_group_bin_17230 = frame (4k)
frame_vm_group_bin_17231 = frame (4k)
frame_vm_group_bin_17232 = frame (4k)
frame_vm_group_bin_17233 = frame (4k)
frame_vm_group_bin_17234 = frame (4k)
frame_vm_group_bin_17235 = frame (4k)
frame_vm_group_bin_17236 = frame (4k)
frame_vm_group_bin_17237 = frame (4k)
frame_vm_group_bin_17238 = frame (4k)
frame_vm_group_bin_17239 = frame (4k)
frame_vm_group_bin_1724 = frame (4k)
frame_vm_group_bin_17240 = frame (4k)
frame_vm_group_bin_17241 = frame (4k)
frame_vm_group_bin_17242 = frame (4k)
frame_vm_group_bin_17243 = frame (4k)
frame_vm_group_bin_17244 = frame (4k)
frame_vm_group_bin_17245 = frame (4k)
frame_vm_group_bin_17246 = frame (4k)
frame_vm_group_bin_17247 = frame (4k)
frame_vm_group_bin_17248 = frame (4k)
frame_vm_group_bin_17249 = frame (4k)
frame_vm_group_bin_1725 = frame (4k)
frame_vm_group_bin_17250 = frame (4k)
frame_vm_group_bin_17251 = frame (4k)
frame_vm_group_bin_17252 = frame (4k)
frame_vm_group_bin_17253 = frame (4k)
frame_vm_group_bin_17254 = frame (4k)
frame_vm_group_bin_17255 = frame (4k)
frame_vm_group_bin_17256 = frame (4k)
frame_vm_group_bin_17257 = frame (4k)
frame_vm_group_bin_17258 = frame (4k)
frame_vm_group_bin_17259 = frame (4k)
frame_vm_group_bin_1726 = frame (4k)
frame_vm_group_bin_17260 = frame (4k)
frame_vm_group_bin_17261 = frame (4k)
frame_vm_group_bin_17262 = frame (4k)
frame_vm_group_bin_17263 = frame (4k)
frame_vm_group_bin_17264 = frame (4k)
frame_vm_group_bin_17265 = frame (4k)
frame_vm_group_bin_17266 = frame (4k)
frame_vm_group_bin_17267 = frame (4k)
frame_vm_group_bin_17268 = frame (4k)
frame_vm_group_bin_17269 = frame (4k)
frame_vm_group_bin_1727 = frame (4k)
frame_vm_group_bin_17270 = frame (4k)
frame_vm_group_bin_17271 = frame (4k)
frame_vm_group_bin_17272 = frame (4k)
frame_vm_group_bin_17273 = frame (4k)
frame_vm_group_bin_17274 = frame (4k)
frame_vm_group_bin_17275 = frame (4k)
frame_vm_group_bin_17276 = frame (4k)
frame_vm_group_bin_17277 = frame (4k)
frame_vm_group_bin_17278 = frame (4k)
frame_vm_group_bin_17279 = frame (4k)
frame_vm_group_bin_1728 = frame (4k)
frame_vm_group_bin_17280 = frame (4k)
frame_vm_group_bin_17281 = frame (4k)
frame_vm_group_bin_17282 = frame (4k)
frame_vm_group_bin_17283 = frame (4k)
frame_vm_group_bin_17284 = frame (4k)
frame_vm_group_bin_17285 = frame (4k)
frame_vm_group_bin_17286 = frame (4k)
frame_vm_group_bin_17287 = frame (4k)
frame_vm_group_bin_17288 = frame (4k)
frame_vm_group_bin_17289 = frame (4k)
frame_vm_group_bin_1729 = frame (4k)
frame_vm_group_bin_17290 = frame (4k)
frame_vm_group_bin_17291 = frame (4k)
frame_vm_group_bin_17292 = frame (4k)
frame_vm_group_bin_17293 = frame (4k)
frame_vm_group_bin_17294 = frame (4k)
frame_vm_group_bin_17295 = frame (4k)
frame_vm_group_bin_17296 = frame (4k)
frame_vm_group_bin_17297 = frame (4k)
frame_vm_group_bin_17298 = frame (4k)
frame_vm_group_bin_17299 = frame (4k)
frame_vm_group_bin_1730 = frame (4k)
frame_vm_group_bin_17300 = frame (4k)
frame_vm_group_bin_17301 = frame (4k)
frame_vm_group_bin_17302 = frame (4k)
frame_vm_group_bin_17303 = frame (4k)
frame_vm_group_bin_17304 = frame (4k)
frame_vm_group_bin_17305 = frame (4k)
frame_vm_group_bin_17306 = frame (4k)
frame_vm_group_bin_17307 = frame (4k)
frame_vm_group_bin_17308 = frame (4k)
frame_vm_group_bin_17309 = frame (4k)
frame_vm_group_bin_1731 = frame (4k)
frame_vm_group_bin_17310 = frame (4k)
frame_vm_group_bin_17311 = frame (4k)
frame_vm_group_bin_17312 = frame (4k)
frame_vm_group_bin_17313 = frame (4k)
frame_vm_group_bin_17314 = frame (4k)
frame_vm_group_bin_17315 = frame (4k)
frame_vm_group_bin_17316 = frame (4k)
frame_vm_group_bin_17317 = frame (4k)
frame_vm_group_bin_17318 = frame (4k)
frame_vm_group_bin_17319 = frame (4k)
frame_vm_group_bin_1732 = frame (4k)
frame_vm_group_bin_17320 = frame (4k)
frame_vm_group_bin_17321 = frame (4k)
frame_vm_group_bin_17322 = frame (4k)
frame_vm_group_bin_17323 = frame (4k)
frame_vm_group_bin_17324 = frame (4k)
frame_vm_group_bin_17325 = frame (4k)
frame_vm_group_bin_17326 = frame (4k)
frame_vm_group_bin_17327 = frame (4k)
frame_vm_group_bin_17328 = frame (4k)
frame_vm_group_bin_17329 = frame (4k)
frame_vm_group_bin_1733 = frame (4k)
frame_vm_group_bin_17330 = frame (4k)
frame_vm_group_bin_17331 = frame (4k)
frame_vm_group_bin_17332 = frame (4k)
frame_vm_group_bin_17333 = frame (4k)
frame_vm_group_bin_17334 = frame (4k)
frame_vm_group_bin_17335 = frame (4k)
frame_vm_group_bin_17336 = frame (4k)
frame_vm_group_bin_17337 = frame (4k)
frame_vm_group_bin_17338 = frame (4k)
frame_vm_group_bin_17339 = frame (4k)
frame_vm_group_bin_1734 = frame (4k)
frame_vm_group_bin_17340 = frame (4k)
frame_vm_group_bin_17341 = frame (4k)
frame_vm_group_bin_17342 = frame (4k)
frame_vm_group_bin_17343 = frame (4k)
frame_vm_group_bin_17344 = frame (4k)
frame_vm_group_bin_17345 = frame (4k)
frame_vm_group_bin_17346 = frame (4k)
frame_vm_group_bin_17347 = frame (4k)
frame_vm_group_bin_17348 = frame (4k)
frame_vm_group_bin_17349 = frame (4k)
frame_vm_group_bin_1735 = frame (4k)
frame_vm_group_bin_17350 = frame (4k)
frame_vm_group_bin_17351 = frame (4k)
frame_vm_group_bin_17352 = frame (4k)
frame_vm_group_bin_17353 = frame (4k)
frame_vm_group_bin_17354 = frame (4k)
frame_vm_group_bin_17355 = frame (4k)
frame_vm_group_bin_17356 = frame (4k)
frame_vm_group_bin_17357 = frame (4k)
frame_vm_group_bin_17358 = frame (4k)
frame_vm_group_bin_17359 = frame (4k)
frame_vm_group_bin_1736 = frame (4k)
frame_vm_group_bin_17360 = frame (4k)
frame_vm_group_bin_17361 = frame (4k)
frame_vm_group_bin_17362 = frame (4k)
frame_vm_group_bin_17363 = frame (4k)
frame_vm_group_bin_17364 = frame (4k)
frame_vm_group_bin_17365 = frame (4k)
frame_vm_group_bin_17366 = frame (4k)
frame_vm_group_bin_17367 = frame (4k)
frame_vm_group_bin_17368 = frame (4k)
frame_vm_group_bin_17369 = frame (4k)
frame_vm_group_bin_1737 = frame (4k)
frame_vm_group_bin_17370 = frame (4k)
frame_vm_group_bin_17371 = frame (4k)
frame_vm_group_bin_17372 = frame (4k)
frame_vm_group_bin_17373 = frame (4k)
frame_vm_group_bin_17374 = frame (4k)
frame_vm_group_bin_17375 = frame (4k)
frame_vm_group_bin_17376 = frame (4k)
frame_vm_group_bin_17377 = frame (4k)
frame_vm_group_bin_17378 = frame (4k)
frame_vm_group_bin_17379 = frame (4k)
frame_vm_group_bin_1738 = frame (4k)
frame_vm_group_bin_17380 = frame (4k)
frame_vm_group_bin_17381 = frame (4k)
frame_vm_group_bin_17382 = frame (4k)
frame_vm_group_bin_17383 = frame (4k)
frame_vm_group_bin_17384 = frame (4k)
frame_vm_group_bin_17385 = frame (4k)
frame_vm_group_bin_17386 = frame (4k)
frame_vm_group_bin_17387 = frame (4k)
frame_vm_group_bin_17388 = frame (4k)
frame_vm_group_bin_17389 = frame (4k)
frame_vm_group_bin_1739 = frame (4k)
frame_vm_group_bin_17390 = frame (4k)
frame_vm_group_bin_17391 = frame (4k)
frame_vm_group_bin_17392 = frame (4k)
frame_vm_group_bin_17393 = frame (4k)
frame_vm_group_bin_17394 = frame (4k)
frame_vm_group_bin_17395 = frame (4k)
frame_vm_group_bin_17396 = frame (4k)
frame_vm_group_bin_17397 = frame (4k)
frame_vm_group_bin_17398 = frame (4k)
frame_vm_group_bin_17399 = frame (4k)
frame_vm_group_bin_1740 = frame (4k)
frame_vm_group_bin_17400 = frame (4k)
frame_vm_group_bin_17401 = frame (4k)
frame_vm_group_bin_17402 = frame (4k)
frame_vm_group_bin_17403 = frame (4k)
frame_vm_group_bin_17404 = frame (4k)
frame_vm_group_bin_17405 = frame (4k)
frame_vm_group_bin_17406 = frame (4k)
frame_vm_group_bin_17407 = frame (4k)
frame_vm_group_bin_17408 = frame (4k)
frame_vm_group_bin_17409 = frame (4k)
frame_vm_group_bin_1741 = frame (4k)
frame_vm_group_bin_17410 = frame (4k)
frame_vm_group_bin_17411 = frame (4k)
frame_vm_group_bin_17412 = frame (4k)
frame_vm_group_bin_17413 = frame (4k)
frame_vm_group_bin_17414 = frame (4k)
frame_vm_group_bin_17415 = frame (4k)
frame_vm_group_bin_17416 = frame (4k)
frame_vm_group_bin_17417 = frame (4k)
frame_vm_group_bin_17418 = frame (4k)
frame_vm_group_bin_17419 = frame (4k)
frame_vm_group_bin_1742 = frame (4k)
frame_vm_group_bin_17420 = frame (4k)
frame_vm_group_bin_17421 = frame (4k)
frame_vm_group_bin_17422 = frame (4k)
frame_vm_group_bin_17423 = frame (4k)
frame_vm_group_bin_17424 = frame (4k)
frame_vm_group_bin_17425 = frame (4k)
frame_vm_group_bin_17426 = frame (4k)
frame_vm_group_bin_17427 = frame (4k)
frame_vm_group_bin_17428 = frame (4k)
frame_vm_group_bin_17429 = frame (4k)
frame_vm_group_bin_1743 = frame (4k)
frame_vm_group_bin_17430 = frame (4k)
frame_vm_group_bin_17431 = frame (4k)
frame_vm_group_bin_17432 = frame (4k)
frame_vm_group_bin_17433 = frame (4k)
frame_vm_group_bin_17434 = frame (4k)
frame_vm_group_bin_17435 = frame (4k)
frame_vm_group_bin_17436 = frame (4k)
frame_vm_group_bin_17437 = frame (4k)
frame_vm_group_bin_17438 = frame (4k)
frame_vm_group_bin_17439 = frame (4k)
frame_vm_group_bin_1744 = frame (4k)
frame_vm_group_bin_17440 = frame (4k)
frame_vm_group_bin_17441 = frame (4k)
frame_vm_group_bin_17442 = frame (4k)
frame_vm_group_bin_17443 = frame (4k)
frame_vm_group_bin_17444 = frame (4k)
frame_vm_group_bin_17445 = frame (4k)
frame_vm_group_bin_17446 = frame (4k)
frame_vm_group_bin_17447 = frame (4k)
frame_vm_group_bin_17448 = frame (4k)
frame_vm_group_bin_17449 = frame (4k)
frame_vm_group_bin_1745 = frame (4k)
frame_vm_group_bin_17450 = frame (4k)
frame_vm_group_bin_17451 = frame (4k)
frame_vm_group_bin_17452 = frame (4k)
frame_vm_group_bin_17453 = frame (4k)
frame_vm_group_bin_17454 = frame (4k)
frame_vm_group_bin_17455 = frame (4k)
frame_vm_group_bin_17456 = frame (4k)
frame_vm_group_bin_17457 = frame (4k)
frame_vm_group_bin_17458 = frame (4k)
frame_vm_group_bin_17459 = frame (4k)
frame_vm_group_bin_1746 = frame (4k)
frame_vm_group_bin_17460 = frame (4k)
frame_vm_group_bin_17461 = frame (4k)
frame_vm_group_bin_17462 = frame (4k)
frame_vm_group_bin_17463 = frame (4k)
frame_vm_group_bin_17464 = frame (4k)
frame_vm_group_bin_17465 = frame (4k)
frame_vm_group_bin_17466 = frame (4k)
frame_vm_group_bin_17467 = frame (4k)
frame_vm_group_bin_17468 = frame (4k)
frame_vm_group_bin_17469 = frame (4k)
frame_vm_group_bin_1747 = frame (4k)
frame_vm_group_bin_17470 = frame (4k)
frame_vm_group_bin_17471 = frame (4k)
frame_vm_group_bin_17472 = frame (4k)
frame_vm_group_bin_17473 = frame (4k)
frame_vm_group_bin_17474 = frame (4k)
frame_vm_group_bin_17475 = frame (4k)
frame_vm_group_bin_17476 = frame (4k)
frame_vm_group_bin_17477 = frame (4k)
frame_vm_group_bin_17478 = frame (4k)
frame_vm_group_bin_17479 = frame (4k)
frame_vm_group_bin_1748 = frame (4k)
frame_vm_group_bin_17480 = frame (4k)
frame_vm_group_bin_17481 = frame (4k)
frame_vm_group_bin_17482 = frame (4k)
frame_vm_group_bin_17483 = frame (4k)
frame_vm_group_bin_17484 = frame (4k)
frame_vm_group_bin_17485 = frame (4k)
frame_vm_group_bin_17486 = frame (4k)
frame_vm_group_bin_17487 = frame (4k)
frame_vm_group_bin_17488 = frame (4k)
frame_vm_group_bin_17489 = frame (4k)
frame_vm_group_bin_1749 = frame (4k)
frame_vm_group_bin_17490 = frame (4k)
frame_vm_group_bin_17491 = frame (4k)
frame_vm_group_bin_17492 = frame (4k)
frame_vm_group_bin_17493 = frame (4k)
frame_vm_group_bin_17494 = frame (4k)
frame_vm_group_bin_17495 = frame (4k)
frame_vm_group_bin_17496 = frame (4k)
frame_vm_group_bin_17497 = frame (4k)
frame_vm_group_bin_17498 = frame (4k)
frame_vm_group_bin_17499 = frame (4k)
frame_vm_group_bin_1750 = frame (4k)
frame_vm_group_bin_17500 = frame (4k)
frame_vm_group_bin_17501 = frame (4k)
frame_vm_group_bin_17502 = frame (4k)
frame_vm_group_bin_17503 = frame (4k)
frame_vm_group_bin_17504 = frame (4k)
frame_vm_group_bin_17505 = frame (4k)
frame_vm_group_bin_17506 = frame (4k)
frame_vm_group_bin_17507 = frame (4k)
frame_vm_group_bin_17508 = frame (4k)
frame_vm_group_bin_17509 = frame (4k)
frame_vm_group_bin_1751 = frame (4k)
frame_vm_group_bin_17510 = frame (4k)
frame_vm_group_bin_17511 = frame (4k)
frame_vm_group_bin_17512 = frame (4k)
frame_vm_group_bin_17513 = frame (4k)
frame_vm_group_bin_17514 = frame (4k)
frame_vm_group_bin_17515 = frame (4k)
frame_vm_group_bin_17516 = frame (4k)
frame_vm_group_bin_17517 = frame (4k)
frame_vm_group_bin_17518 = frame (4k)
frame_vm_group_bin_17519 = frame (4k)
frame_vm_group_bin_1752 = frame (4k)
frame_vm_group_bin_17520 = frame (4k)
frame_vm_group_bin_17521 = frame (4k)
frame_vm_group_bin_17522 = frame (4k)
frame_vm_group_bin_17523 = frame (4k)
frame_vm_group_bin_17524 = frame (4k)
frame_vm_group_bin_17525 = frame (4k)
frame_vm_group_bin_17526 = frame (4k)
frame_vm_group_bin_17527 = frame (4k)
frame_vm_group_bin_17528 = frame (4k)
frame_vm_group_bin_17529 = frame (4k)
frame_vm_group_bin_1753 = frame (4k)
frame_vm_group_bin_17530 = frame (4k)
frame_vm_group_bin_17531 = frame (4k)
frame_vm_group_bin_17532 = frame (4k)
frame_vm_group_bin_17533 = frame (4k)
frame_vm_group_bin_17534 = frame (4k)
frame_vm_group_bin_17535 = frame (4k)
frame_vm_group_bin_17536 = frame (4k)
frame_vm_group_bin_17537 = frame (4k)
frame_vm_group_bin_17538 = frame (4k)
frame_vm_group_bin_17539 = frame (4k)
frame_vm_group_bin_1754 = frame (4k)
frame_vm_group_bin_17540 = frame (4k)
frame_vm_group_bin_17541 = frame (4k)
frame_vm_group_bin_17542 = frame (4k)
frame_vm_group_bin_17543 = frame (4k)
frame_vm_group_bin_17544 = frame (4k)
frame_vm_group_bin_17545 = frame (4k)
frame_vm_group_bin_17546 = frame (4k)
frame_vm_group_bin_17547 = frame (4k)
frame_vm_group_bin_17548 = frame (4k)
frame_vm_group_bin_17549 = frame (4k)
frame_vm_group_bin_1755 = frame (4k)
frame_vm_group_bin_17550 = frame (4k)
frame_vm_group_bin_17551 = frame (4k)
frame_vm_group_bin_17552 = frame (4k)
frame_vm_group_bin_17553 = frame (4k)
frame_vm_group_bin_17554 = frame (4k)
frame_vm_group_bin_17555 = frame (4k)
frame_vm_group_bin_17556 = frame (4k)
frame_vm_group_bin_17557 = frame (4k)
frame_vm_group_bin_17558 = frame (4k)
frame_vm_group_bin_17559 = frame (4k)
frame_vm_group_bin_1756 = frame (4k)
frame_vm_group_bin_17560 = frame (4k)
frame_vm_group_bin_17561 = frame (4k)
frame_vm_group_bin_17562 = frame (4k)
frame_vm_group_bin_17563 = frame (4k)
frame_vm_group_bin_17564 = frame (4k)
frame_vm_group_bin_17565 = frame (4k)
frame_vm_group_bin_17566 = frame (4k)
frame_vm_group_bin_17567 = frame (4k)
frame_vm_group_bin_17568 = frame (4k)
frame_vm_group_bin_17569 = frame (4k)
frame_vm_group_bin_1757 = frame (4k)
frame_vm_group_bin_17570 = frame (4k)
frame_vm_group_bin_17571 = frame (4k)
frame_vm_group_bin_17572 = frame (4k)
frame_vm_group_bin_17573 = frame (4k)
frame_vm_group_bin_17574 = frame (4k)
frame_vm_group_bin_17575 = frame (4k)
frame_vm_group_bin_17576 = frame (4k)
frame_vm_group_bin_17577 = frame (4k)
frame_vm_group_bin_17578 = frame (4k)
frame_vm_group_bin_17579 = frame (4k)
frame_vm_group_bin_1758 = frame (4k)
frame_vm_group_bin_17580 = frame (4k)
frame_vm_group_bin_17581 = frame (4k)
frame_vm_group_bin_17582 = frame (4k)
frame_vm_group_bin_17583 = frame (4k)
frame_vm_group_bin_17584 = frame (4k)
frame_vm_group_bin_17585 = frame (4k)
frame_vm_group_bin_17586 = frame (4k)
frame_vm_group_bin_17587 = frame (4k)
frame_vm_group_bin_17588 = frame (4k)
frame_vm_group_bin_17589 = frame (4k)
frame_vm_group_bin_1759 = frame (4k)
frame_vm_group_bin_17590 = frame (4k)
frame_vm_group_bin_17591 = frame (4k)
frame_vm_group_bin_17592 = frame (4k)
frame_vm_group_bin_17593 = frame (4k)
frame_vm_group_bin_17594 = frame (4k)
frame_vm_group_bin_17595 = frame (4k)
frame_vm_group_bin_17596 = frame (4k)
frame_vm_group_bin_17597 = frame (4k)
frame_vm_group_bin_17598 = frame (4k)
frame_vm_group_bin_17599 = frame (4k)
frame_vm_group_bin_1760 = frame (4k)
frame_vm_group_bin_17600 = frame (4k)
frame_vm_group_bin_17601 = frame (4k)
frame_vm_group_bin_17602 = frame (4k)
frame_vm_group_bin_17603 = frame (4k)
frame_vm_group_bin_17604 = frame (4k)
frame_vm_group_bin_17605 = frame (4k)
frame_vm_group_bin_17606 = frame (4k)
frame_vm_group_bin_17607 = frame (4k)
frame_vm_group_bin_17608 = frame (4k)
frame_vm_group_bin_17609 = frame (4k)
frame_vm_group_bin_1761 = frame (4k)
frame_vm_group_bin_17610 = frame (4k)
frame_vm_group_bin_17611 = frame (4k)
frame_vm_group_bin_17612 = frame (4k)
frame_vm_group_bin_17613 = frame (4k)
frame_vm_group_bin_17614 = frame (4k)
frame_vm_group_bin_17615 = frame (4k)
frame_vm_group_bin_17616 = frame (4k)
frame_vm_group_bin_17617 = frame (4k)
frame_vm_group_bin_17618 = frame (4k)
frame_vm_group_bin_17619 = frame (4k)
frame_vm_group_bin_1762 = frame (4k)
frame_vm_group_bin_17620 = frame (4k)
frame_vm_group_bin_17621 = frame (4k)
frame_vm_group_bin_17622 = frame (4k)
frame_vm_group_bin_17623 = frame (4k)
frame_vm_group_bin_17624 = frame (4k)
frame_vm_group_bin_17625 = frame (4k)
frame_vm_group_bin_17626 = frame (4k)
frame_vm_group_bin_17627 = frame (4k)
frame_vm_group_bin_17628 = frame (4k)
frame_vm_group_bin_17629 = frame (4k)
frame_vm_group_bin_1763 = frame (4k)
frame_vm_group_bin_17630 = frame (4k)
frame_vm_group_bin_17631 = frame (4k)
frame_vm_group_bin_17632 = frame (4k)
frame_vm_group_bin_17633 = frame (4k)
frame_vm_group_bin_17634 = frame (4k)
frame_vm_group_bin_17635 = frame (4k)
frame_vm_group_bin_17636 = frame (4k)
frame_vm_group_bin_17637 = frame (4k)
frame_vm_group_bin_17638 = frame (4k)
frame_vm_group_bin_17639 = frame (4k)
frame_vm_group_bin_1764 = frame (4k)
frame_vm_group_bin_17640 = frame (4k)
frame_vm_group_bin_17641 = frame (4k)
frame_vm_group_bin_17642 = frame (4k)
frame_vm_group_bin_17643 = frame (4k)
frame_vm_group_bin_17644 = frame (4k)
frame_vm_group_bin_17645 = frame (4k)
frame_vm_group_bin_17646 = frame (4k)
frame_vm_group_bin_17647 = frame (4k)
frame_vm_group_bin_17648 = frame (4k)
frame_vm_group_bin_17649 = frame (4k)
frame_vm_group_bin_1765 = frame (4k)
frame_vm_group_bin_17650 = frame (4k)
frame_vm_group_bin_17651 = frame (4k)
frame_vm_group_bin_17652 = frame (4k)
frame_vm_group_bin_17653 = frame (4k)
frame_vm_group_bin_17654 = frame (4k)
frame_vm_group_bin_17655 = frame (4k)
frame_vm_group_bin_17656 = frame (4k)
frame_vm_group_bin_17657 = frame (4k)
frame_vm_group_bin_17658 = frame (4k)
frame_vm_group_bin_17659 = frame (4k)
frame_vm_group_bin_1766 = frame (4k)
frame_vm_group_bin_17660 = frame (4k)
frame_vm_group_bin_17661 = frame (4k)
frame_vm_group_bin_17662 = frame (4k)
frame_vm_group_bin_17663 = frame (4k)
frame_vm_group_bin_17664 = frame (4k)
frame_vm_group_bin_17665 = frame (4k)
frame_vm_group_bin_17666 = frame (4k)
frame_vm_group_bin_17667 = frame (4k)
frame_vm_group_bin_17668 = frame (4k)
frame_vm_group_bin_17669 = frame (4k)
frame_vm_group_bin_1767 = frame (4k)
frame_vm_group_bin_17670 = frame (4k)
frame_vm_group_bin_17671 = frame (4k)
frame_vm_group_bin_17672 = frame (4k)
frame_vm_group_bin_17673 = frame (4k)
frame_vm_group_bin_17674 = frame (4k)
frame_vm_group_bin_17675 = frame (4k)
frame_vm_group_bin_17676 = frame (4k)
frame_vm_group_bin_17677 = frame (4k)
frame_vm_group_bin_17678 = frame (4k)
frame_vm_group_bin_17679 = frame (4k)
frame_vm_group_bin_1768 = frame (4k)
frame_vm_group_bin_17680 = frame (4k)
frame_vm_group_bin_17681 = frame (4k)
frame_vm_group_bin_17682 = frame (4k)
frame_vm_group_bin_17683 = frame (4k)
frame_vm_group_bin_17684 = frame (4k)
frame_vm_group_bin_17685 = frame (4k)
frame_vm_group_bin_17686 = frame (4k)
frame_vm_group_bin_17687 = frame (4k)
frame_vm_group_bin_17688 = frame (4k)
frame_vm_group_bin_17689 = frame (4k)
frame_vm_group_bin_1769 = frame (4k)
frame_vm_group_bin_17690 = frame (4k)
frame_vm_group_bin_17691 = frame (4k)
frame_vm_group_bin_17692 = frame (4k)
frame_vm_group_bin_17693 = frame (4k)
frame_vm_group_bin_17694 = frame (4k)
frame_vm_group_bin_17695 = frame (4k)
frame_vm_group_bin_17696 = frame (4k)
frame_vm_group_bin_17697 = frame (4k)
frame_vm_group_bin_17698 = frame (4k)
frame_vm_group_bin_17699 = frame (4k)
frame_vm_group_bin_1770 = frame (4k)
frame_vm_group_bin_17700 = frame (4k)
frame_vm_group_bin_17701 = frame (4k)
frame_vm_group_bin_17702 = frame (4k)
frame_vm_group_bin_17703 = frame (4k)
frame_vm_group_bin_17704 = frame (4k)
frame_vm_group_bin_17705 = frame (4k)
frame_vm_group_bin_17706 = frame (4k)
frame_vm_group_bin_17707 = frame (4k)
frame_vm_group_bin_17708 = frame (4k)
frame_vm_group_bin_17709 = frame (4k)
frame_vm_group_bin_1771 = frame (4k)
frame_vm_group_bin_17710 = frame (4k)
frame_vm_group_bin_17711 = frame (4k)
frame_vm_group_bin_17712 = frame (4k)
frame_vm_group_bin_17713 = frame (4k)
frame_vm_group_bin_17714 = frame (4k)
frame_vm_group_bin_17715 = frame (4k)
frame_vm_group_bin_17716 = frame (4k)
frame_vm_group_bin_17717 = frame (4k)
frame_vm_group_bin_17718 = frame (4k)
frame_vm_group_bin_17719 = frame (4k)
frame_vm_group_bin_1772 = frame (4k)
frame_vm_group_bin_17720 = frame (4k)
frame_vm_group_bin_17721 = frame (4k)
frame_vm_group_bin_17722 = frame (4k)
frame_vm_group_bin_17723 = frame (4k)
frame_vm_group_bin_17724 = frame (4k)
frame_vm_group_bin_17725 = frame (4k)
frame_vm_group_bin_17726 = frame (4k)
frame_vm_group_bin_17727 = frame (4k)
frame_vm_group_bin_17728 = frame (4k)
frame_vm_group_bin_17729 = frame (4k)
frame_vm_group_bin_1773 = frame (4k)
frame_vm_group_bin_17730 = frame (4k)
frame_vm_group_bin_17731 = frame (4k)
frame_vm_group_bin_17732 = frame (4k)
frame_vm_group_bin_17733 = frame (4k)
frame_vm_group_bin_17734 = frame (4k)
frame_vm_group_bin_17735 = frame (4k)
frame_vm_group_bin_17736 = frame (4k)
frame_vm_group_bin_17737 = frame (4k)
frame_vm_group_bin_17738 = frame (4k)
frame_vm_group_bin_17739 = frame (4k)
frame_vm_group_bin_1774 = frame (4k)
frame_vm_group_bin_17740 = frame (4k)
frame_vm_group_bin_17741 = frame (4k)
frame_vm_group_bin_17742 = frame (4k)
frame_vm_group_bin_17743 = frame (4k)
frame_vm_group_bin_17744 = frame (4k)
frame_vm_group_bin_17745 = frame (4k)
frame_vm_group_bin_17746 = frame (4k)
frame_vm_group_bin_17747 = frame (4k)
frame_vm_group_bin_17748 = frame (4k)
frame_vm_group_bin_17749 = frame (4k)
frame_vm_group_bin_1775 = frame (4k)
frame_vm_group_bin_17750 = frame (4k)
frame_vm_group_bin_17751 = frame (4k)
frame_vm_group_bin_17752 = frame (4k)
frame_vm_group_bin_17753 = frame (4k)
frame_vm_group_bin_17755 = frame (4k)
frame_vm_group_bin_17756 = frame (4k)
frame_vm_group_bin_17757 = frame (4k)
frame_vm_group_bin_17758 = frame (4k)
frame_vm_group_bin_17759 = frame (4k)
frame_vm_group_bin_1776 = frame (4k)
frame_vm_group_bin_17760 = frame (4k)
frame_vm_group_bin_17761 = frame (4k)
frame_vm_group_bin_17762 = frame (4k)
frame_vm_group_bin_17763 = frame (4k)
frame_vm_group_bin_17764 = frame (4k)
frame_vm_group_bin_17765 = frame (4k)
frame_vm_group_bin_17766 = frame (4k)
frame_vm_group_bin_17767 = frame (4k)
frame_vm_group_bin_17768 = frame (4k)
frame_vm_group_bin_17769 = frame (4k)
frame_vm_group_bin_1777 = frame (4k)
frame_vm_group_bin_17770 = frame (4k)
frame_vm_group_bin_17771 = frame (4k)
frame_vm_group_bin_17772 = frame (4k)
frame_vm_group_bin_17773 = frame (4k)
frame_vm_group_bin_17774 = frame (4k)
frame_vm_group_bin_17775 = frame (4k)
frame_vm_group_bin_17776 = frame (4k)
frame_vm_group_bin_17777 = frame (4k)
frame_vm_group_bin_17778 = frame (4k)
frame_vm_group_bin_17779 = frame (4k)
frame_vm_group_bin_1778 = frame (4k)
frame_vm_group_bin_17780 = frame (4k)
frame_vm_group_bin_17781 = frame (4k)
frame_vm_group_bin_17782 = frame (4k)
frame_vm_group_bin_17783 = frame (4k)
frame_vm_group_bin_17784 = frame (4k)
frame_vm_group_bin_17785 = frame (4k)
frame_vm_group_bin_17786 = frame (4k)
frame_vm_group_bin_17787 = frame (4k)
frame_vm_group_bin_17788 = frame (4k)
frame_vm_group_bin_17789 = frame (4k)
frame_vm_group_bin_1779 = frame (4k)
frame_vm_group_bin_17790 = frame (4k)
frame_vm_group_bin_17791 = frame (4k)
frame_vm_group_bin_17792 = frame (4k)
frame_vm_group_bin_17793 = frame (4k)
frame_vm_group_bin_17794 = frame (4k)
frame_vm_group_bin_17795 = frame (4k)
frame_vm_group_bin_17796 = frame (4k)
frame_vm_group_bin_17797 = frame (4k)
frame_vm_group_bin_17798 = frame (4k)
frame_vm_group_bin_17799 = frame (4k)
frame_vm_group_bin_1780 = frame (4k)
frame_vm_group_bin_17800 = frame (4k)
frame_vm_group_bin_17801 = frame (4k)
frame_vm_group_bin_17802 = frame (4k)
frame_vm_group_bin_17803 = frame (4k)
frame_vm_group_bin_17804 = frame (4k)
frame_vm_group_bin_17805 = frame (4k)
frame_vm_group_bin_17806 = frame (4k)
frame_vm_group_bin_17807 = frame (4k)
frame_vm_group_bin_17808 = frame (4k)
frame_vm_group_bin_17809 = frame (4k)
frame_vm_group_bin_1781 = frame (4k)
frame_vm_group_bin_17810 = frame (4k)
frame_vm_group_bin_17811 = frame (4k)
frame_vm_group_bin_17812 = frame (4k)
frame_vm_group_bin_17813 = frame (4k)
frame_vm_group_bin_17814 = frame (4k)
frame_vm_group_bin_17815 = frame (4k)
frame_vm_group_bin_17816 = frame (4k)
frame_vm_group_bin_17817 = frame (4k)
frame_vm_group_bin_17818 = frame (4k)
frame_vm_group_bin_17819 = frame (4k)
frame_vm_group_bin_1782 = frame (4k)
frame_vm_group_bin_17820 = frame (4k)
frame_vm_group_bin_17821 = frame (4k)
frame_vm_group_bin_17822 = frame (4k)
frame_vm_group_bin_17823 = frame (4k)
frame_vm_group_bin_17824 = frame (4k)
frame_vm_group_bin_17825 = frame (4k)
frame_vm_group_bin_17826 = frame (4k)
frame_vm_group_bin_17827 = frame (4k)
frame_vm_group_bin_17828 = frame (4k)
frame_vm_group_bin_17829 = frame (4k)
frame_vm_group_bin_1783 = frame (4k)
frame_vm_group_bin_17830 = frame (4k)
frame_vm_group_bin_17831 = frame (4k)
frame_vm_group_bin_17832 = frame (4k)
frame_vm_group_bin_17833 = frame (4k)
frame_vm_group_bin_17834 = frame (4k)
frame_vm_group_bin_17835 = frame (4k)
frame_vm_group_bin_17836 = frame (4k)
frame_vm_group_bin_17837 = frame (4k)
frame_vm_group_bin_17838 = frame (4k)
frame_vm_group_bin_17839 = frame (4k)
frame_vm_group_bin_1784 = frame (4k)
frame_vm_group_bin_17840 = frame (4k)
frame_vm_group_bin_17841 = frame (4k)
frame_vm_group_bin_17842 = frame (4k)
frame_vm_group_bin_17843 = frame (4k)
frame_vm_group_bin_17844 = frame (4k)
frame_vm_group_bin_17845 = frame (4k)
frame_vm_group_bin_17846 = frame (4k)
frame_vm_group_bin_17847 = frame (4k)
frame_vm_group_bin_17848 = frame (4k)
frame_vm_group_bin_17849 = frame (4k)
frame_vm_group_bin_1785 = frame (4k)
frame_vm_group_bin_17850 = frame (4k)
frame_vm_group_bin_17851 = frame (4k)
frame_vm_group_bin_17852 = frame (4k)
frame_vm_group_bin_17853 = frame (4k)
frame_vm_group_bin_17854 = frame (4k)
frame_vm_group_bin_17855 = frame (4k)
frame_vm_group_bin_17856 = frame (4k)
frame_vm_group_bin_17857 = frame (4k)
frame_vm_group_bin_17858 = frame (4k)
frame_vm_group_bin_17859 = frame (4k)
frame_vm_group_bin_1786 = frame (4k)
frame_vm_group_bin_17860 = frame (4k)
frame_vm_group_bin_17861 = frame (4k)
frame_vm_group_bin_17862 = frame (4k)
frame_vm_group_bin_17863 = frame (4k)
frame_vm_group_bin_17864 = frame (4k)
frame_vm_group_bin_17865 = frame (4k)
frame_vm_group_bin_17866 = frame (4k)
frame_vm_group_bin_17867 = frame (4k)
frame_vm_group_bin_17868 = frame (4k)
frame_vm_group_bin_17869 = frame (4k)
frame_vm_group_bin_1787 = frame (4k)
frame_vm_group_bin_17870 = frame (4k)
frame_vm_group_bin_17871 = frame (4k)
frame_vm_group_bin_17872 = frame (4k)
frame_vm_group_bin_17873 = frame (4k)
frame_vm_group_bin_17874 = frame (4k)
frame_vm_group_bin_17875 = frame (4k)
frame_vm_group_bin_17876 = frame (4k)
frame_vm_group_bin_17877 = frame (4k)
frame_vm_group_bin_17878 = frame (4k)
frame_vm_group_bin_17879 = frame (4k)
frame_vm_group_bin_1788 = frame (4k)
frame_vm_group_bin_17880 = frame (4k)
frame_vm_group_bin_17881 = frame (4k)
frame_vm_group_bin_17882 = frame (4k)
frame_vm_group_bin_17883 = frame (4k)
frame_vm_group_bin_17884 = frame (4k)
frame_vm_group_bin_17885 = frame (4k)
frame_vm_group_bin_17886 = frame (4k)
frame_vm_group_bin_17887 = frame (4k)
frame_vm_group_bin_17888 = frame (4k)
frame_vm_group_bin_17889 = frame (4k)
frame_vm_group_bin_1789 = frame (4k)
frame_vm_group_bin_17890 = frame (4k)
frame_vm_group_bin_17891 = frame (4k)
frame_vm_group_bin_17892 = frame (4k)
frame_vm_group_bin_17893 = frame (4k)
frame_vm_group_bin_17894 = frame (4k)
frame_vm_group_bin_17895 = frame (4k)
frame_vm_group_bin_17896 = frame (4k)
frame_vm_group_bin_17897 = frame (4k)
frame_vm_group_bin_17898 = frame (4k)
frame_vm_group_bin_17899 = frame (4k)
frame_vm_group_bin_1790 = frame (4k)
frame_vm_group_bin_17900 = frame (4k)
frame_vm_group_bin_17901 = frame (4k)
frame_vm_group_bin_17902 = frame (4k)
frame_vm_group_bin_17903 = frame (4k)
frame_vm_group_bin_17904 = frame (4k)
frame_vm_group_bin_17905 = frame (4k)
frame_vm_group_bin_17906 = frame (4k)
frame_vm_group_bin_17907 = frame (4k)
frame_vm_group_bin_17908 = frame (4k)
frame_vm_group_bin_17909 = frame (4k)
frame_vm_group_bin_1791 = frame (4k)
frame_vm_group_bin_17910 = frame (4k)
frame_vm_group_bin_17911 = frame (4k)
frame_vm_group_bin_17912 = frame (4k)
frame_vm_group_bin_17913 = frame (4k)
frame_vm_group_bin_17914 = frame (4k)
frame_vm_group_bin_17915 = frame (4k)
frame_vm_group_bin_17916 = frame (4k)
frame_vm_group_bin_17917 = frame (4k)
frame_vm_group_bin_17918 = frame (4k)
frame_vm_group_bin_17919 = frame (4k)
frame_vm_group_bin_1792 = frame (4k)
frame_vm_group_bin_17920 = frame (4k)
frame_vm_group_bin_17921 = frame (4k)
frame_vm_group_bin_17922 = frame (4k)
frame_vm_group_bin_17923 = frame (4k)
frame_vm_group_bin_17924 = frame (4k)
frame_vm_group_bin_17925 = frame (4k)
frame_vm_group_bin_17926 = frame (4k)
frame_vm_group_bin_17927 = frame (4k)
frame_vm_group_bin_17928 = frame (4k)
frame_vm_group_bin_17929 = frame (4k)
frame_vm_group_bin_1793 = frame (4k)
frame_vm_group_bin_17930 = frame (4k)
frame_vm_group_bin_17931 = frame (4k)
frame_vm_group_bin_17932 = frame (4k)
frame_vm_group_bin_17933 = frame (4k)
frame_vm_group_bin_17934 = frame (4k)
frame_vm_group_bin_17935 = frame (4k)
frame_vm_group_bin_17936 = frame (4k)
frame_vm_group_bin_17937 = frame (4k)
frame_vm_group_bin_17938 = frame (4k)
frame_vm_group_bin_17939 = frame (4k)
frame_vm_group_bin_1794 = frame (4k)
frame_vm_group_bin_17940 = frame (4k)
frame_vm_group_bin_17941 = frame (4k)
frame_vm_group_bin_17942 = frame (4k)
frame_vm_group_bin_17943 = frame (4k)
frame_vm_group_bin_17944 = frame (4k)
frame_vm_group_bin_17945 = frame (4k)
frame_vm_group_bin_17946 = frame (4k)
frame_vm_group_bin_17947 = frame (4k)
frame_vm_group_bin_17948 = frame (4k)
frame_vm_group_bin_17949 = frame (4k)
frame_vm_group_bin_1795 = frame (4k)
frame_vm_group_bin_17950 = frame (4k)
frame_vm_group_bin_17951 = frame (4k)
frame_vm_group_bin_17952 = frame (4k)
frame_vm_group_bin_17953 = frame (4k)
frame_vm_group_bin_17954 = frame (4k)
frame_vm_group_bin_17955 = frame (4k)
frame_vm_group_bin_17956 = frame (4k)
frame_vm_group_bin_17957 = frame (4k)
frame_vm_group_bin_17958 = frame (4k)
frame_vm_group_bin_17959 = frame (4k)
frame_vm_group_bin_1796 = frame (4k)
frame_vm_group_bin_17960 = frame (4k)
frame_vm_group_bin_17961 = frame (4k)
frame_vm_group_bin_17962 = frame (4k)
frame_vm_group_bin_17963 = frame (4k)
frame_vm_group_bin_17964 = frame (4k)
frame_vm_group_bin_17965 = frame (4k)
frame_vm_group_bin_17966 = frame (4k)
frame_vm_group_bin_17967 = frame (4k)
frame_vm_group_bin_17968 = frame (4k)
frame_vm_group_bin_17969 = frame (4k)
frame_vm_group_bin_1797 = frame (4k)
frame_vm_group_bin_17970 = frame (4k)
frame_vm_group_bin_17971 = frame (4k)
frame_vm_group_bin_17972 = frame (4k)
frame_vm_group_bin_17973 = frame (4k)
frame_vm_group_bin_17974 = frame (4k)
frame_vm_group_bin_17975 = frame (4k)
frame_vm_group_bin_17976 = frame (4k)
frame_vm_group_bin_17977 = frame (4k)
frame_vm_group_bin_17978 = frame (4k)
frame_vm_group_bin_17979 = frame (4k)
frame_vm_group_bin_1798 = frame (4k)
frame_vm_group_bin_17980 = frame (4k)
frame_vm_group_bin_17981 = frame (4k)
frame_vm_group_bin_17982 = frame (4k)
frame_vm_group_bin_17983 = frame (4k)
frame_vm_group_bin_17984 = frame (4k)
frame_vm_group_bin_17985 = frame (4k)
frame_vm_group_bin_17986 = frame (4k)
frame_vm_group_bin_17987 = frame (4k)
frame_vm_group_bin_17988 = frame (4k)
frame_vm_group_bin_17989 = frame (4k)
frame_vm_group_bin_1799 = frame (4k)
frame_vm_group_bin_17990 = frame (4k)
frame_vm_group_bin_17991 = frame (4k)
frame_vm_group_bin_17992 = frame (4k)
frame_vm_group_bin_17993 = frame (4k)
frame_vm_group_bin_17994 = frame (4k)
frame_vm_group_bin_17995 = frame (4k)
frame_vm_group_bin_17996 = frame (4k)
frame_vm_group_bin_17997 = frame (4k)
frame_vm_group_bin_17998 = frame (4k)
frame_vm_group_bin_17999 = frame (4k)
frame_vm_group_bin_1800 = frame (4k)
frame_vm_group_bin_18000 = frame (4k)
frame_vm_group_bin_18001 = frame (4k)
frame_vm_group_bin_18002 = frame (4k)
frame_vm_group_bin_18003 = frame (4k)
frame_vm_group_bin_18004 = frame (4k)
frame_vm_group_bin_18005 = frame (4k)
frame_vm_group_bin_18006 = frame (4k)
frame_vm_group_bin_18007 = frame (4k)
frame_vm_group_bin_18008 = frame (4k)
frame_vm_group_bin_18009 = frame (4k)
frame_vm_group_bin_1801 = frame (4k)
frame_vm_group_bin_18010 = frame (4k)
frame_vm_group_bin_18011 = frame (4k)
frame_vm_group_bin_18012 = frame (4k)
frame_vm_group_bin_18013 = frame (4k)
frame_vm_group_bin_18014 = frame (4k)
frame_vm_group_bin_18015 = frame (4k)
frame_vm_group_bin_18016 = frame (4k)
frame_vm_group_bin_18017 = frame (4k)
frame_vm_group_bin_18018 = frame (4k)
frame_vm_group_bin_18019 = frame (4k)
frame_vm_group_bin_1802 = frame (4k)
frame_vm_group_bin_18020 = frame (4k)
frame_vm_group_bin_18021 = frame (4k)
frame_vm_group_bin_18022 = frame (4k)
frame_vm_group_bin_18023 = frame (4k)
frame_vm_group_bin_18024 = frame (4k)
frame_vm_group_bin_18025 = frame (4k)
frame_vm_group_bin_18026 = frame (4k)
frame_vm_group_bin_18027 = frame (4k)
frame_vm_group_bin_18028 = frame (4k)
frame_vm_group_bin_18029 = frame (4k)
frame_vm_group_bin_1803 = frame (4k)
frame_vm_group_bin_18030 = frame (4k)
frame_vm_group_bin_18031 = frame (4k)
frame_vm_group_bin_18032 = frame (4k)
frame_vm_group_bin_18033 = frame (4k)
frame_vm_group_bin_18034 = frame (4k)
frame_vm_group_bin_18035 = frame (4k)
frame_vm_group_bin_18036 = frame (4k)
frame_vm_group_bin_18037 = frame (4k)
frame_vm_group_bin_18038 = frame (4k)
frame_vm_group_bin_18039 = frame (4k)
frame_vm_group_bin_1804 = frame (4k)
frame_vm_group_bin_18040 = frame (4k)
frame_vm_group_bin_18041 = frame (4k)
frame_vm_group_bin_18042 = frame (4k)
frame_vm_group_bin_18043 = frame (4k)
frame_vm_group_bin_18044 = frame (4k)
frame_vm_group_bin_18045 = frame (4k)
frame_vm_group_bin_18046 = frame (4k)
frame_vm_group_bin_18047 = frame (4k)
frame_vm_group_bin_18048 = frame (4k)
frame_vm_group_bin_18049 = frame (4k)
frame_vm_group_bin_1805 = frame (4k)
frame_vm_group_bin_18050 = frame (4k)
frame_vm_group_bin_18051 = frame (4k)
frame_vm_group_bin_18052 = frame (4k)
frame_vm_group_bin_18053 = frame (4k)
frame_vm_group_bin_18054 = frame (4k)
frame_vm_group_bin_18055 = frame (4k)
frame_vm_group_bin_18056 = frame (4k)
frame_vm_group_bin_18057 = frame (4k)
frame_vm_group_bin_18058 = frame (4k)
frame_vm_group_bin_18059 = frame (4k)
frame_vm_group_bin_1806 = frame (4k)
frame_vm_group_bin_18060 = frame (4k)
frame_vm_group_bin_18061 = frame (4k)
frame_vm_group_bin_18062 = frame (4k)
frame_vm_group_bin_18063 = frame (4k)
frame_vm_group_bin_18064 = frame (4k)
frame_vm_group_bin_18065 = frame (4k)
frame_vm_group_bin_18066 = frame (4k)
frame_vm_group_bin_18067 = frame (4k)
frame_vm_group_bin_18068 = frame (4k)
frame_vm_group_bin_18069 = frame (4k)
frame_vm_group_bin_1807 = frame (4k)
frame_vm_group_bin_18070 = frame (4k)
frame_vm_group_bin_18071 = frame (4k)
frame_vm_group_bin_18072 = frame (4k)
frame_vm_group_bin_18073 = frame (4k)
frame_vm_group_bin_18074 = frame (4k)
frame_vm_group_bin_18075 = frame (4k)
frame_vm_group_bin_18076 = frame (4k)
frame_vm_group_bin_18077 = frame (4k)
frame_vm_group_bin_18078 = frame (4k)
frame_vm_group_bin_18079 = frame (4k)
frame_vm_group_bin_1808 = frame (4k)
frame_vm_group_bin_18080 = frame (4k)
frame_vm_group_bin_18081 = frame (4k)
frame_vm_group_bin_18082 = frame (4k)
frame_vm_group_bin_18083 = frame (4k)
frame_vm_group_bin_18084 = frame (4k)
frame_vm_group_bin_18085 = frame (4k)
frame_vm_group_bin_18086 = frame (4k)
frame_vm_group_bin_18087 = frame (4k)
frame_vm_group_bin_18088 = frame (4k)
frame_vm_group_bin_18089 = frame (4k)
frame_vm_group_bin_1809 = frame (4k)
frame_vm_group_bin_18090 = frame (4k)
frame_vm_group_bin_18091 = frame (4k)
frame_vm_group_bin_18092 = frame (4k)
frame_vm_group_bin_18093 = frame (4k)
frame_vm_group_bin_18094 = frame (4k)
frame_vm_group_bin_18095 = frame (4k)
frame_vm_group_bin_18096 = frame (4k)
frame_vm_group_bin_18097 = frame (4k)
frame_vm_group_bin_18098 = frame (4k)
frame_vm_group_bin_18099 = frame (4k)
frame_vm_group_bin_1810 = frame (4k)
frame_vm_group_bin_18100 = frame (4k)
frame_vm_group_bin_18101 = frame (4k)
frame_vm_group_bin_18102 = frame (4k)
frame_vm_group_bin_18103 = frame (4k)
frame_vm_group_bin_18104 = frame (4k)
frame_vm_group_bin_18105 = frame (4k)
frame_vm_group_bin_18106 = frame (4k)
frame_vm_group_bin_18107 = frame (4k)
frame_vm_group_bin_18108 = frame (4k)
frame_vm_group_bin_18109 = frame (4k)
frame_vm_group_bin_1811 = frame (4k)
frame_vm_group_bin_18110 = frame (4k)
frame_vm_group_bin_18111 = frame (4k)
frame_vm_group_bin_18112 = frame (4k)
frame_vm_group_bin_18113 = frame (4k)
frame_vm_group_bin_18114 = frame (4k)
frame_vm_group_bin_18115 = frame (4k)
frame_vm_group_bin_18116 = frame (4k)
frame_vm_group_bin_18117 = frame (4k)
frame_vm_group_bin_18118 = frame (4k)
frame_vm_group_bin_18119 = frame (4k)
frame_vm_group_bin_1812 = frame (4k)
frame_vm_group_bin_18120 = frame (4k)
frame_vm_group_bin_18121 = frame (4k)
frame_vm_group_bin_18122 = frame (4k)
frame_vm_group_bin_18123 = frame (4k)
frame_vm_group_bin_18124 = frame (4k)
frame_vm_group_bin_18125 = frame (4k)
frame_vm_group_bin_18126 = frame (4k)
frame_vm_group_bin_18127 = frame (4k)
frame_vm_group_bin_18128 = frame (4k)
frame_vm_group_bin_18129 = frame (4k)
frame_vm_group_bin_1813 = frame (4k)
frame_vm_group_bin_18130 = frame (4k)
frame_vm_group_bin_18131 = frame (4k)
frame_vm_group_bin_18132 = frame (4k)
frame_vm_group_bin_18133 = frame (4k)
frame_vm_group_bin_18134 = frame (4k)
frame_vm_group_bin_18135 = frame (4k)
frame_vm_group_bin_18136 = frame (4k)
frame_vm_group_bin_18137 = frame (4k)
frame_vm_group_bin_18138 = frame (4k)
frame_vm_group_bin_18139 = frame (4k)
frame_vm_group_bin_1814 = frame (4k)
frame_vm_group_bin_18140 = frame (4k)
frame_vm_group_bin_18141 = frame (4k)
frame_vm_group_bin_18142 = frame (4k)
frame_vm_group_bin_18143 = frame (4k)
frame_vm_group_bin_18144 = frame (4k)
frame_vm_group_bin_18145 = frame (4k)
frame_vm_group_bin_18146 = frame (4k)
frame_vm_group_bin_18147 = frame (4k)
frame_vm_group_bin_18148 = frame (4k)
frame_vm_group_bin_18149 = frame (4k)
frame_vm_group_bin_1815 = frame (4k)
frame_vm_group_bin_18150 = frame (4k)
frame_vm_group_bin_18151 = frame (4k)
frame_vm_group_bin_18152 = frame (4k)
frame_vm_group_bin_18153 = frame (4k)
frame_vm_group_bin_18154 = frame (4k)
frame_vm_group_bin_18155 = frame (4k)
frame_vm_group_bin_18156 = frame (4k)
frame_vm_group_bin_18157 = frame (4k)
frame_vm_group_bin_18158 = frame (4k)
frame_vm_group_bin_18159 = frame (4k)
frame_vm_group_bin_1816 = frame (4k)
frame_vm_group_bin_18160 = frame (4k)
frame_vm_group_bin_18161 = frame (4k)
frame_vm_group_bin_18162 = frame (4k)
frame_vm_group_bin_18163 = frame (4k)
frame_vm_group_bin_18164 = frame (4k)
frame_vm_group_bin_18165 = frame (4k)
frame_vm_group_bin_18166 = frame (4k)
frame_vm_group_bin_18167 = frame (4k)
frame_vm_group_bin_18168 = frame (4k)
frame_vm_group_bin_18169 = frame (4k)
frame_vm_group_bin_1817 = frame (4k)
frame_vm_group_bin_18170 = frame (4k)
frame_vm_group_bin_18171 = frame (4k)
frame_vm_group_bin_18172 = frame (4k)
frame_vm_group_bin_18173 = frame (4k)
frame_vm_group_bin_18174 = frame (4k)
frame_vm_group_bin_18175 = frame (4k)
frame_vm_group_bin_18176 = frame (4k)
frame_vm_group_bin_18177 = frame (4k)
frame_vm_group_bin_18178 = frame (4k)
frame_vm_group_bin_18179 = frame (4k)
frame_vm_group_bin_1818 = frame (4k)
frame_vm_group_bin_18180 = frame (4k)
frame_vm_group_bin_18181 = frame (4k)
frame_vm_group_bin_18182 = frame (4k)
frame_vm_group_bin_18183 = frame (4k)
frame_vm_group_bin_18184 = frame (4k)
frame_vm_group_bin_18185 = frame (4k)
frame_vm_group_bin_18186 = frame (4k)
frame_vm_group_bin_18187 = frame (4k)
frame_vm_group_bin_18188 = frame (4k)
frame_vm_group_bin_18189 = frame (4k)
frame_vm_group_bin_1819 = frame (4k)
frame_vm_group_bin_18190 = frame (4k)
frame_vm_group_bin_18191 = frame (4k)
frame_vm_group_bin_18192 = frame (4k)
frame_vm_group_bin_18193 = frame (4k)
frame_vm_group_bin_18194 = frame (4k)
frame_vm_group_bin_18195 = frame (4k)
frame_vm_group_bin_18196 = frame (4k)
frame_vm_group_bin_18197 = frame (4k)
frame_vm_group_bin_18198 = frame (4k)
frame_vm_group_bin_18199 = frame (4k)
frame_vm_group_bin_1820 = frame (4k)
frame_vm_group_bin_18200 = frame (4k)
frame_vm_group_bin_18201 = frame (4k)
frame_vm_group_bin_18202 = frame (4k)
frame_vm_group_bin_18203 = frame (4k)
frame_vm_group_bin_18204 = frame (4k)
frame_vm_group_bin_18205 = frame (4k)
frame_vm_group_bin_18206 = frame (4k)
frame_vm_group_bin_18207 = frame (4k)
frame_vm_group_bin_18208 = frame (4k)
frame_vm_group_bin_18209 = frame (4k)
frame_vm_group_bin_1821 = frame (4k)
frame_vm_group_bin_18210 = frame (4k)
frame_vm_group_bin_18211 = frame (4k)
frame_vm_group_bin_18212 = frame (4k)
frame_vm_group_bin_18213 = frame (4k)
frame_vm_group_bin_18214 = frame (4k)
frame_vm_group_bin_18215 = frame (4k)
frame_vm_group_bin_18216 = frame (4k)
frame_vm_group_bin_18217 = frame (4k)
frame_vm_group_bin_18218 = frame (4k)
frame_vm_group_bin_18219 = frame (4k)
frame_vm_group_bin_1822 = frame (4k)
frame_vm_group_bin_18220 = frame (4k)
frame_vm_group_bin_18221 = frame (4k)
frame_vm_group_bin_18222 = frame (4k)
frame_vm_group_bin_18223 = frame (4k)
frame_vm_group_bin_18224 = frame (4k)
frame_vm_group_bin_18225 = frame (4k)
frame_vm_group_bin_18226 = frame (4k)
frame_vm_group_bin_18227 = frame (4k)
frame_vm_group_bin_18228 = frame (4k)
frame_vm_group_bin_18229 = frame (4k)
frame_vm_group_bin_1823 = frame (4k)
frame_vm_group_bin_18230 = frame (4k)
frame_vm_group_bin_18231 = frame (4k)
frame_vm_group_bin_18232 = frame (4k)
frame_vm_group_bin_18233 = frame (4k)
frame_vm_group_bin_18234 = frame (4k)
frame_vm_group_bin_18235 = frame (4k)
frame_vm_group_bin_18236 = frame (4k)
frame_vm_group_bin_18237 = frame (4k)
frame_vm_group_bin_18238 = frame (4k)
frame_vm_group_bin_18239 = frame (4k)
frame_vm_group_bin_1824 = frame (4k)
frame_vm_group_bin_18240 = frame (4k)
frame_vm_group_bin_18241 = frame (4k)
frame_vm_group_bin_18242 = frame (4k)
frame_vm_group_bin_18243 = frame (4k)
frame_vm_group_bin_18244 = frame (4k)
frame_vm_group_bin_18245 = frame (4k)
frame_vm_group_bin_18246 = frame (4k)
frame_vm_group_bin_18247 = frame (4k)
frame_vm_group_bin_18248 = frame (4k)
frame_vm_group_bin_18249 = frame (4k)
frame_vm_group_bin_1825 = frame (4k)
frame_vm_group_bin_18250 = frame (4k)
frame_vm_group_bin_18251 = frame (4k)
frame_vm_group_bin_18252 = frame (4k)
frame_vm_group_bin_18253 = frame (4k)
frame_vm_group_bin_18254 = frame (4k)
frame_vm_group_bin_18255 = frame (4k)
frame_vm_group_bin_18256 = frame (4k)
frame_vm_group_bin_18257 = frame (4k)
frame_vm_group_bin_18258 = frame (4k)
frame_vm_group_bin_18259 = frame (4k)
frame_vm_group_bin_1826 = frame (4k)
frame_vm_group_bin_18260 = frame (4k)
frame_vm_group_bin_18261 = frame (4k)
frame_vm_group_bin_18262 = frame (4k)
frame_vm_group_bin_18263 = frame (4k)
frame_vm_group_bin_18264 = frame (4k)
frame_vm_group_bin_18265 = frame (4k)
frame_vm_group_bin_18266 = frame (4k)
frame_vm_group_bin_18267 = frame (4k)
frame_vm_group_bin_18268 = frame (4k)
frame_vm_group_bin_18269 = frame (4k)
frame_vm_group_bin_1827 = frame (4k)
frame_vm_group_bin_18270 = frame (4k)
frame_vm_group_bin_18271 = frame (4k)
frame_vm_group_bin_18272 = frame (4k)
frame_vm_group_bin_18273 = frame (4k)
frame_vm_group_bin_18274 = frame (4k)
frame_vm_group_bin_18275 = frame (4k)
frame_vm_group_bin_18276 = frame (4k)
frame_vm_group_bin_18277 = frame (4k)
frame_vm_group_bin_18278 = frame (4k)
frame_vm_group_bin_18279 = frame (4k)
frame_vm_group_bin_1828 = frame (4k)
frame_vm_group_bin_18280 = frame (4k)
frame_vm_group_bin_18281 = frame (4k)
frame_vm_group_bin_18282 = frame (4k)
frame_vm_group_bin_18283 = frame (4k)
frame_vm_group_bin_18284 = frame (4k)
frame_vm_group_bin_18285 = frame (4k)
frame_vm_group_bin_18286 = frame (4k)
frame_vm_group_bin_18287 = frame (4k)
frame_vm_group_bin_18288 = frame (4k)
frame_vm_group_bin_18289 = frame (4k)
frame_vm_group_bin_1829 = frame (4k)
frame_vm_group_bin_18290 = frame (4k)
frame_vm_group_bin_18291 = frame (4k)
frame_vm_group_bin_18292 = frame (4k)
frame_vm_group_bin_18293 = frame (4k)
frame_vm_group_bin_18294 = frame (4k)
frame_vm_group_bin_18295 = frame (4k)
frame_vm_group_bin_18296 = frame (4k)
frame_vm_group_bin_18297 = frame (4k)
frame_vm_group_bin_18298 = frame (4k)
frame_vm_group_bin_18299 = frame (4k)
frame_vm_group_bin_1830 = frame (4k)
frame_vm_group_bin_18300 = frame (4k)
frame_vm_group_bin_18301 = frame (4k)
frame_vm_group_bin_18302 = frame (4k)
frame_vm_group_bin_18303 = frame (4k)
frame_vm_group_bin_18304 = frame (4k)
frame_vm_group_bin_18305 = frame (4k)
frame_vm_group_bin_18306 = frame (4k)
frame_vm_group_bin_18307 = frame (4k)
frame_vm_group_bin_18308 = frame (4k)
frame_vm_group_bin_18309 = frame (4k)
frame_vm_group_bin_1831 = frame (4k)
frame_vm_group_bin_18310 = frame (4k)
frame_vm_group_bin_18311 = frame (4k)
frame_vm_group_bin_18312 = frame (4k)
frame_vm_group_bin_18313 = frame (4k)
frame_vm_group_bin_18314 = frame (4k)
frame_vm_group_bin_18315 = frame (4k)
frame_vm_group_bin_18316 = frame (4k)
frame_vm_group_bin_18317 = frame (4k)
frame_vm_group_bin_18318 = frame (4k)
frame_vm_group_bin_18319 = frame (4k)
frame_vm_group_bin_1832 = frame (4k)
frame_vm_group_bin_18320 = frame (4k)
frame_vm_group_bin_18321 = frame (4k)
frame_vm_group_bin_18322 = frame (4k)
frame_vm_group_bin_18323 = frame (4k)
frame_vm_group_bin_18324 = frame (4k)
frame_vm_group_bin_18325 = frame (4k)
frame_vm_group_bin_18326 = frame (4k)
frame_vm_group_bin_18327 = frame (4k)
frame_vm_group_bin_18328 = frame (4k)
frame_vm_group_bin_18329 = frame (4k)
frame_vm_group_bin_1833 = frame (4k)
frame_vm_group_bin_18330 = frame (4k)
frame_vm_group_bin_18331 = frame (4k)
frame_vm_group_bin_18332 = frame (4k)
frame_vm_group_bin_18333 = frame (4k)
frame_vm_group_bin_18334 = frame (4k)
frame_vm_group_bin_18335 = frame (4k)
frame_vm_group_bin_18336 = frame (4k)
frame_vm_group_bin_18337 = frame (4k)
frame_vm_group_bin_18338 = frame (4k)
frame_vm_group_bin_18339 = frame (4k)
frame_vm_group_bin_1834 = frame (4k)
frame_vm_group_bin_18340 = frame (4k)
frame_vm_group_bin_18341 = frame (4k)
frame_vm_group_bin_18342 = frame (4k)
frame_vm_group_bin_18343 = frame (4k)
frame_vm_group_bin_18344 = frame (4k)
frame_vm_group_bin_18345 = frame (4k)
frame_vm_group_bin_18346 = frame (4k)
frame_vm_group_bin_18347 = frame (4k)
frame_vm_group_bin_18348 = frame (4k)
frame_vm_group_bin_18349 = frame (4k)
frame_vm_group_bin_1835 = frame (4k)
frame_vm_group_bin_18350 = frame (4k)
frame_vm_group_bin_18351 = frame (4k)
frame_vm_group_bin_18352 = frame (4k)
frame_vm_group_bin_18353 = frame (4k)
frame_vm_group_bin_18354 = frame (4k)
frame_vm_group_bin_18355 = frame (4k)
frame_vm_group_bin_18356 = frame (4k)
frame_vm_group_bin_18357 = frame (4k)
frame_vm_group_bin_18358 = frame (4k)
frame_vm_group_bin_18359 = frame (4k)
frame_vm_group_bin_1836 = frame (4k)
frame_vm_group_bin_18360 = frame (4k)
frame_vm_group_bin_18361 = frame (4k)
frame_vm_group_bin_18362 = frame (4k)
frame_vm_group_bin_18363 = frame (4k)
frame_vm_group_bin_18364 = frame (4k)
frame_vm_group_bin_18365 = frame (4k)
frame_vm_group_bin_18366 = frame (4k)
frame_vm_group_bin_18367 = frame (4k)
frame_vm_group_bin_18368 = frame (4k)
frame_vm_group_bin_18369 = frame (4k)
frame_vm_group_bin_1837 = frame (4k)
frame_vm_group_bin_18370 = frame (4k)
frame_vm_group_bin_18371 = frame (4k)
frame_vm_group_bin_18372 = frame (4k)
frame_vm_group_bin_18373 = frame (4k)
frame_vm_group_bin_18374 = frame (4k)
frame_vm_group_bin_18375 = frame (4k)
frame_vm_group_bin_18376 = frame (4k)
frame_vm_group_bin_18377 = frame (4k)
frame_vm_group_bin_18378 = frame (4k)
frame_vm_group_bin_18379 = frame (4k)
frame_vm_group_bin_1838 = frame (4k)
frame_vm_group_bin_18380 = frame (4k)
frame_vm_group_bin_18381 = frame (4k)
frame_vm_group_bin_18382 = frame (4k)
frame_vm_group_bin_18383 = frame (4k)
frame_vm_group_bin_18384 = frame (4k)
frame_vm_group_bin_18385 = frame (4k)
frame_vm_group_bin_18386 = frame (4k)
frame_vm_group_bin_18387 = frame (4k)
frame_vm_group_bin_18388 = frame (4k)
frame_vm_group_bin_18389 = frame (4k)
frame_vm_group_bin_1839 = frame (4k)
frame_vm_group_bin_18390 = frame (4k)
frame_vm_group_bin_18391 = frame (4k)
frame_vm_group_bin_18392 = frame (4k)
frame_vm_group_bin_18393 = frame (4k)
frame_vm_group_bin_18394 = frame (4k)
frame_vm_group_bin_18395 = frame (4k)
frame_vm_group_bin_18396 = frame (4k)
frame_vm_group_bin_18397 = frame (4k)
frame_vm_group_bin_18398 = frame (4k)
frame_vm_group_bin_18399 = frame (4k)
frame_vm_group_bin_1840 = frame (4k)
frame_vm_group_bin_18400 = frame (4k)
frame_vm_group_bin_18401 = frame (4k)
frame_vm_group_bin_18402 = frame (4k)
frame_vm_group_bin_18403 = frame (4k)
frame_vm_group_bin_18404 = frame (4k)
frame_vm_group_bin_18405 = frame (4k)
frame_vm_group_bin_18406 = frame (4k)
frame_vm_group_bin_18407 = frame (4k)
frame_vm_group_bin_18408 = frame (4k)
frame_vm_group_bin_18409 = frame (4k)
frame_vm_group_bin_1841 = frame (4k)
frame_vm_group_bin_18410 = frame (4k)
frame_vm_group_bin_18411 = frame (4k)
frame_vm_group_bin_18412 = frame (4k)
frame_vm_group_bin_18413 = frame (4k)
frame_vm_group_bin_18414 = frame (4k)
frame_vm_group_bin_18415 = frame (4k)
frame_vm_group_bin_18416 = frame (4k)
frame_vm_group_bin_18417 = frame (4k)
frame_vm_group_bin_18418 = frame (4k)
frame_vm_group_bin_18419 = frame (4k)
frame_vm_group_bin_1842 = frame (4k)
frame_vm_group_bin_18420 = frame (4k)
frame_vm_group_bin_18421 = frame (4k)
frame_vm_group_bin_18422 = frame (4k)
frame_vm_group_bin_18423 = frame (4k)
frame_vm_group_bin_18424 = frame (4k)
frame_vm_group_bin_18425 = frame (4k)
frame_vm_group_bin_18426 = frame (4k)
frame_vm_group_bin_18427 = frame (4k)
frame_vm_group_bin_18428 = frame (4k)
frame_vm_group_bin_18429 = frame (4k)
frame_vm_group_bin_1843 = frame (4k)
frame_vm_group_bin_18430 = frame (4k)
frame_vm_group_bin_18431 = frame (4k)
frame_vm_group_bin_18432 = frame (4k)
frame_vm_group_bin_18433 = frame (4k)
frame_vm_group_bin_18434 = frame (4k)
frame_vm_group_bin_18435 = frame (4k)
frame_vm_group_bin_18436 = frame (4k)
frame_vm_group_bin_18437 = frame (4k)
frame_vm_group_bin_18438 = frame (4k)
frame_vm_group_bin_18439 = frame (4k)
frame_vm_group_bin_1844 = frame (4k)
frame_vm_group_bin_18440 = frame (4k)
frame_vm_group_bin_18441 = frame (4k)
frame_vm_group_bin_18442 = frame (4k)
frame_vm_group_bin_18443 = frame (4k)
frame_vm_group_bin_18444 = frame (4k)
frame_vm_group_bin_18445 = frame (4k)
frame_vm_group_bin_18446 = frame (4k)
frame_vm_group_bin_18447 = frame (4k)
frame_vm_group_bin_18448 = frame (4k)
frame_vm_group_bin_18449 = frame (4k)
frame_vm_group_bin_1845 = frame (4k)
frame_vm_group_bin_18450 = frame (4k)
frame_vm_group_bin_18451 = frame (4k)
frame_vm_group_bin_18452 = frame (4k)
frame_vm_group_bin_18453 = frame (4k)
frame_vm_group_bin_18454 = frame (4k)
frame_vm_group_bin_18455 = frame (4k)
frame_vm_group_bin_18456 = frame (4k)
frame_vm_group_bin_18457 = frame (4k)
frame_vm_group_bin_18458 = frame (4k)
frame_vm_group_bin_18459 = frame (4k)
frame_vm_group_bin_1846 = frame (4k)
frame_vm_group_bin_18460 = frame (4k)
frame_vm_group_bin_18461 = frame (4k)
frame_vm_group_bin_18462 = frame (4k)
frame_vm_group_bin_18463 = frame (4k)
frame_vm_group_bin_18464 = frame (4k)
frame_vm_group_bin_18465 = frame (4k)
frame_vm_group_bin_18466 = frame (4k)
frame_vm_group_bin_18467 = frame (4k)
frame_vm_group_bin_18468 = frame (4k)
frame_vm_group_bin_18469 = frame (4k)
frame_vm_group_bin_1847 = frame (4k)
frame_vm_group_bin_18470 = frame (4k)
frame_vm_group_bin_18471 = frame (4k)
frame_vm_group_bin_18472 = frame (4k)
frame_vm_group_bin_18473 = frame (4k)
frame_vm_group_bin_18474 = frame (4k)
frame_vm_group_bin_18475 = frame (4k)
frame_vm_group_bin_18476 = frame (4k)
frame_vm_group_bin_18477 = frame (4k)
frame_vm_group_bin_18478 = frame (4k)
frame_vm_group_bin_18479 = frame (4k)
frame_vm_group_bin_1848 = frame (4k)
frame_vm_group_bin_18480 = frame (4k)
frame_vm_group_bin_18481 = frame (4k)
frame_vm_group_bin_18482 = frame (4k)
frame_vm_group_bin_18483 = frame (4k)
frame_vm_group_bin_18484 = frame (4k)
frame_vm_group_bin_18485 = frame (4k)
frame_vm_group_bin_18486 = frame (4k)
frame_vm_group_bin_18487 = frame (4k)
frame_vm_group_bin_18488 = frame (4k)
frame_vm_group_bin_18489 = frame (4k)
frame_vm_group_bin_1849 = frame (4k)
frame_vm_group_bin_18490 = frame (4k)
frame_vm_group_bin_18491 = frame (4k)
frame_vm_group_bin_18492 = frame (4k)
frame_vm_group_bin_18493 = frame (4k)
frame_vm_group_bin_18494 = frame (4k)
frame_vm_group_bin_18495 = frame (4k)
frame_vm_group_bin_18496 = frame (4k)
frame_vm_group_bin_18497 = frame (4k)
frame_vm_group_bin_18498 = frame (4k)
frame_vm_group_bin_18499 = frame (4k)
frame_vm_group_bin_1850 = frame (4k)
frame_vm_group_bin_18500 = frame (4k)
frame_vm_group_bin_18501 = frame (4k)
frame_vm_group_bin_18502 = frame (4k)
frame_vm_group_bin_18503 = frame (4k)
frame_vm_group_bin_18504 = frame (4k)
frame_vm_group_bin_18505 = frame (4k)
frame_vm_group_bin_18506 = frame (4k)
frame_vm_group_bin_18507 = frame (4k)
frame_vm_group_bin_18508 = frame (4k)
frame_vm_group_bin_18509 = frame (4k)
frame_vm_group_bin_1851 = frame (4k)
frame_vm_group_bin_18510 = frame (4k)
frame_vm_group_bin_18511 = frame (4k)
frame_vm_group_bin_18512 = frame (4k)
frame_vm_group_bin_18513 = frame (4k)
frame_vm_group_bin_18514 = frame (4k)
frame_vm_group_bin_18515 = frame (4k)
frame_vm_group_bin_18516 = frame (4k)
frame_vm_group_bin_18517 = frame (4k)
frame_vm_group_bin_18518 = frame (4k)
frame_vm_group_bin_18519 = frame (4k)
frame_vm_group_bin_1852 = frame (4k)
frame_vm_group_bin_18520 = frame (4k)
frame_vm_group_bin_18521 = frame (4k)
frame_vm_group_bin_18522 = frame (4k)
frame_vm_group_bin_18523 = frame (4k)
frame_vm_group_bin_18524 = frame (4k)
frame_vm_group_bin_18525 = frame (4k)
frame_vm_group_bin_18526 = frame (4k)
frame_vm_group_bin_18527 = frame (4k)
frame_vm_group_bin_18528 = frame (4k)
frame_vm_group_bin_18529 = frame (4k)
frame_vm_group_bin_1853 = frame (4k)
frame_vm_group_bin_18530 = frame (4k)
frame_vm_group_bin_18531 = frame (4k)
frame_vm_group_bin_18532 = frame (4k)
frame_vm_group_bin_18533 = frame (4k)
frame_vm_group_bin_18534 = frame (4k)
frame_vm_group_bin_18535 = frame (4k)
frame_vm_group_bin_18536 = frame (4k)
frame_vm_group_bin_18537 = frame (4k)
frame_vm_group_bin_18538 = frame (4k)
frame_vm_group_bin_18539 = frame (4k)
frame_vm_group_bin_1854 = frame (4k)
frame_vm_group_bin_18540 = frame (4k)
frame_vm_group_bin_18541 = frame (4k)
frame_vm_group_bin_18542 = frame (4k)
frame_vm_group_bin_18543 = frame (4k)
frame_vm_group_bin_18544 = frame (4k)
frame_vm_group_bin_18545 = frame (4k)
frame_vm_group_bin_18546 = frame (4k)
frame_vm_group_bin_18547 = frame (4k)
frame_vm_group_bin_18548 = frame (4k)
frame_vm_group_bin_18549 = frame (4k)
frame_vm_group_bin_1855 = frame (4k)
frame_vm_group_bin_18550 = frame (4k)
frame_vm_group_bin_18551 = frame (4k)
frame_vm_group_bin_18552 = frame (4k)
frame_vm_group_bin_18553 = frame (4k)
frame_vm_group_bin_18554 = frame (4k)
frame_vm_group_bin_18555 = frame (4k)
frame_vm_group_bin_18556 = frame (4k)
frame_vm_group_bin_18557 = frame (4k)
frame_vm_group_bin_18558 = frame (4k)
frame_vm_group_bin_18559 = frame (4k)
frame_vm_group_bin_1856 = frame (4k)
frame_vm_group_bin_18560 = frame (4k)
frame_vm_group_bin_18561 = frame (4k)
frame_vm_group_bin_18562 = frame (4k)
frame_vm_group_bin_18563 = frame (4k)
frame_vm_group_bin_18564 = frame (4k)
frame_vm_group_bin_18565 = frame (4k)
frame_vm_group_bin_18566 = frame (4k)
frame_vm_group_bin_18567 = frame (4k)
frame_vm_group_bin_18568 = frame (4k)
frame_vm_group_bin_18569 = frame (4k)
frame_vm_group_bin_1857 = frame (4k)
frame_vm_group_bin_18570 = frame (4k)
frame_vm_group_bin_18571 = frame (4k)
frame_vm_group_bin_18572 = frame (4k)
frame_vm_group_bin_18573 = frame (4k)
frame_vm_group_bin_18574 = frame (4k)
frame_vm_group_bin_18575 = frame (4k)
frame_vm_group_bin_18576 = frame (4k)
frame_vm_group_bin_18577 = frame (4k)
frame_vm_group_bin_18578 = frame (4k)
frame_vm_group_bin_18579 = frame (4k)
frame_vm_group_bin_1858 = frame (4k)
frame_vm_group_bin_18580 = frame (4k)
frame_vm_group_bin_18581 = frame (4k)
frame_vm_group_bin_18582 = frame (4k)
frame_vm_group_bin_18583 = frame (4k)
frame_vm_group_bin_18584 = frame (4k)
frame_vm_group_bin_18585 = frame (4k)
frame_vm_group_bin_18586 = frame (4k)
frame_vm_group_bin_18587 = frame (4k)
frame_vm_group_bin_18588 = frame (4k)
frame_vm_group_bin_18589 = frame (4k)
frame_vm_group_bin_1859 = frame (4k)
frame_vm_group_bin_18590 = frame (4k)
frame_vm_group_bin_18591 = frame (4k)
frame_vm_group_bin_18592 = frame (4k)
frame_vm_group_bin_18593 = frame (4k)
frame_vm_group_bin_18594 = frame (4k)
frame_vm_group_bin_18595 = frame (4k)
frame_vm_group_bin_18596 = frame (4k)
frame_vm_group_bin_18597 = frame (4k)
frame_vm_group_bin_18598 = frame (4k)
frame_vm_group_bin_18599 = frame (4k)
frame_vm_group_bin_1860 = frame (4k)
frame_vm_group_bin_18600 = frame (4k)
frame_vm_group_bin_18601 = frame (4k)
frame_vm_group_bin_18602 = frame (4k)
frame_vm_group_bin_18603 = frame (4k)
frame_vm_group_bin_18604 = frame (4k)
frame_vm_group_bin_18605 = frame (4k)
frame_vm_group_bin_18606 = frame (4k)
frame_vm_group_bin_18607 = frame (4k)
frame_vm_group_bin_18608 = frame (4k)
frame_vm_group_bin_18609 = frame (4k)
frame_vm_group_bin_1861 = frame (4k)
frame_vm_group_bin_18610 = frame (4k)
frame_vm_group_bin_18611 = frame (4k)
frame_vm_group_bin_18612 = frame (4k)
frame_vm_group_bin_18613 = frame (4k)
frame_vm_group_bin_18614 = frame (4k)
frame_vm_group_bin_18615 = frame (4k)
frame_vm_group_bin_18616 = frame (4k)
frame_vm_group_bin_18617 = frame (4k)
frame_vm_group_bin_18618 = frame (4k)
frame_vm_group_bin_18619 = frame (4k)
frame_vm_group_bin_1862 = frame (4k)
frame_vm_group_bin_18620 = frame (4k)
frame_vm_group_bin_18621 = frame (4k)
frame_vm_group_bin_18622 = frame (4k)
frame_vm_group_bin_18623 = frame (4k)
frame_vm_group_bin_18624 = frame (4k)
frame_vm_group_bin_18625 = frame (4k)
frame_vm_group_bin_18626 = frame (4k)
frame_vm_group_bin_18627 = frame (4k)
frame_vm_group_bin_18628 = frame (4k)
frame_vm_group_bin_18629 = frame (4k)
frame_vm_group_bin_1863 = frame (4k)
frame_vm_group_bin_18630 = frame (4k)
frame_vm_group_bin_18631 = frame (4k)
frame_vm_group_bin_18632 = frame (4k)
frame_vm_group_bin_18633 = frame (4k)
frame_vm_group_bin_18634 = frame (4k)
frame_vm_group_bin_18635 = frame (4k)
frame_vm_group_bin_18636 = frame (4k)
frame_vm_group_bin_18637 = frame (4k)
frame_vm_group_bin_18638 = frame (4k)
frame_vm_group_bin_18639 = frame (4k)
frame_vm_group_bin_1864 = frame (4k)
frame_vm_group_bin_18640 = frame (4k)
frame_vm_group_bin_18641 = frame (4k)
frame_vm_group_bin_18642 = frame (4k)
frame_vm_group_bin_18643 = frame (4k)
frame_vm_group_bin_18644 = frame (4k)
frame_vm_group_bin_18645 = frame (4k)
frame_vm_group_bin_18646 = frame (4k)
frame_vm_group_bin_18647 = frame (4k)
frame_vm_group_bin_18648 = frame (4k)
frame_vm_group_bin_18649 = frame (4k)
frame_vm_group_bin_1865 = frame (4k)
frame_vm_group_bin_18650 = frame (4k)
frame_vm_group_bin_18651 = frame (4k)
frame_vm_group_bin_18652 = frame (4k)
frame_vm_group_bin_18653 = frame (4k)
frame_vm_group_bin_18654 = frame (4k)
frame_vm_group_bin_18655 = frame (4k)
frame_vm_group_bin_18656 = frame (4k)
frame_vm_group_bin_18657 = frame (4k)
frame_vm_group_bin_18658 = frame (4k)
frame_vm_group_bin_18659 = frame (4k)
frame_vm_group_bin_1866 = frame (4k)
frame_vm_group_bin_18660 = frame (4k)
frame_vm_group_bin_18661 = frame (4k)
frame_vm_group_bin_18662 = frame (4k)
frame_vm_group_bin_18663 = frame (4k)
frame_vm_group_bin_18664 = frame (4k)
frame_vm_group_bin_18665 = frame (4k)
frame_vm_group_bin_18666 = frame (4k)
frame_vm_group_bin_18667 = frame (4k)
frame_vm_group_bin_18668 = frame (4k)
frame_vm_group_bin_18669 = frame (4k)
frame_vm_group_bin_1867 = frame (4k)
frame_vm_group_bin_18670 = frame (4k)
frame_vm_group_bin_18671 = frame (4k)
frame_vm_group_bin_18672 = frame (4k)
frame_vm_group_bin_18673 = frame (4k)
frame_vm_group_bin_18674 = frame (4k)
frame_vm_group_bin_18675 = frame (4k)
frame_vm_group_bin_18676 = frame (4k)
frame_vm_group_bin_18677 = frame (4k)
frame_vm_group_bin_18678 = frame (4k)
frame_vm_group_bin_18679 = frame (4k)
frame_vm_group_bin_1868 = frame (4k)
frame_vm_group_bin_18680 = frame (4k)
frame_vm_group_bin_18681 = frame (4k)
frame_vm_group_bin_18682 = frame (4k)
frame_vm_group_bin_18683 = frame (4k)
frame_vm_group_bin_18684 = frame (4k)
frame_vm_group_bin_18685 = frame (4k)
frame_vm_group_bin_18686 = frame (4k)
frame_vm_group_bin_18687 = frame (4k)
frame_vm_group_bin_18688 = frame (4k)
frame_vm_group_bin_18689 = frame (4k)
frame_vm_group_bin_1869 = frame (4k)
frame_vm_group_bin_18690 = frame (4k)
frame_vm_group_bin_18691 = frame (4k)
frame_vm_group_bin_18692 = frame (4k)
frame_vm_group_bin_18693 = frame (4k)
frame_vm_group_bin_18694 = frame (4k)
frame_vm_group_bin_18695 = frame (4k)
frame_vm_group_bin_18696 = frame (4k)
frame_vm_group_bin_18697 = frame (4k)
frame_vm_group_bin_18698 = frame (4k)
frame_vm_group_bin_18699 = frame (4k)
frame_vm_group_bin_1870 = frame (4k)
frame_vm_group_bin_18700 = frame (4k)
frame_vm_group_bin_18701 = frame (4k)
frame_vm_group_bin_18702 = frame (4k)
frame_vm_group_bin_18703 = frame (4k)
frame_vm_group_bin_18704 = frame (4k)
frame_vm_group_bin_18705 = frame (4k)
frame_vm_group_bin_18706 = frame (4k)
frame_vm_group_bin_18707 = frame (4k)
frame_vm_group_bin_18708 = frame (4k)
frame_vm_group_bin_18709 = frame (4k)
frame_vm_group_bin_1871 = frame (4k)
frame_vm_group_bin_18710 = frame (4k)
frame_vm_group_bin_18711 = frame (4k)
frame_vm_group_bin_18712 = frame (4k)
frame_vm_group_bin_18713 = frame (4k)
frame_vm_group_bin_18714 = frame (4k)
frame_vm_group_bin_18715 = frame (4k)
frame_vm_group_bin_18716 = frame (4k)
frame_vm_group_bin_18717 = frame (4k)
frame_vm_group_bin_18718 = frame (4k)
frame_vm_group_bin_18719 = frame (4k)
frame_vm_group_bin_1872 = frame (4k)
frame_vm_group_bin_18720 = frame (4k)
frame_vm_group_bin_18721 = frame (4k)
frame_vm_group_bin_18722 = frame (4k)
frame_vm_group_bin_18723 = frame (4k)
frame_vm_group_bin_18724 = frame (4k)
frame_vm_group_bin_18725 = frame (4k)
frame_vm_group_bin_18726 = frame (4k)
frame_vm_group_bin_18727 = frame (4k)
frame_vm_group_bin_18728 = frame (4k)
frame_vm_group_bin_18729 = frame (4k)
frame_vm_group_bin_1873 = frame (4k)
frame_vm_group_bin_18730 = frame (4k)
frame_vm_group_bin_18731 = frame (4k)
frame_vm_group_bin_18732 = frame (4k)
frame_vm_group_bin_18733 = frame (4k)
frame_vm_group_bin_18734 = frame (4k)
frame_vm_group_bin_18735 = frame (4k)
frame_vm_group_bin_18736 = frame (4k)
frame_vm_group_bin_18737 = frame (4k)
frame_vm_group_bin_18738 = frame (4k)
frame_vm_group_bin_18739 = frame (4k)
frame_vm_group_bin_1874 = frame (4k)
frame_vm_group_bin_18740 = frame (4k)
frame_vm_group_bin_18741 = frame (4k)
frame_vm_group_bin_18742 = frame (4k)
frame_vm_group_bin_18743 = frame (4k)
frame_vm_group_bin_18744 = frame (4k)
frame_vm_group_bin_18745 = frame (4k)
frame_vm_group_bin_18746 = frame (4k)
frame_vm_group_bin_18747 = frame (4k)
frame_vm_group_bin_18748 = frame (4k)
frame_vm_group_bin_18749 = frame (4k)
frame_vm_group_bin_1875 = frame (4k)
frame_vm_group_bin_18750 = frame (4k)
frame_vm_group_bin_18751 = frame (4k)
frame_vm_group_bin_18752 = frame (4k)
frame_vm_group_bin_18753 = frame (4k)
frame_vm_group_bin_18754 = frame (4k)
frame_vm_group_bin_18755 = frame (4k)
frame_vm_group_bin_18756 = frame (4k)
frame_vm_group_bin_18757 = frame (4k)
frame_vm_group_bin_18758 = frame (4k)
frame_vm_group_bin_18759 = frame (4k)
frame_vm_group_bin_1876 = frame (4k)
frame_vm_group_bin_18760 = frame (4k)
frame_vm_group_bin_18761 = frame (4k)
frame_vm_group_bin_18762 = frame (4k)
frame_vm_group_bin_18763 = frame (4k)
frame_vm_group_bin_18764 = frame (4k)
frame_vm_group_bin_18765 = frame (4k)
frame_vm_group_bin_18766 = frame (4k)
frame_vm_group_bin_18767 = frame (4k)
frame_vm_group_bin_18768 = frame (4k)
frame_vm_group_bin_18769 = frame (4k)
frame_vm_group_bin_1877 = frame (4k)
frame_vm_group_bin_18770 = frame (4k)
frame_vm_group_bin_18771 = frame (4k)
frame_vm_group_bin_18772 = frame (4k)
frame_vm_group_bin_18773 = frame (4k)
frame_vm_group_bin_18774 = frame (4k)
frame_vm_group_bin_18775 = frame (4k)
frame_vm_group_bin_18776 = frame (4k)
frame_vm_group_bin_18777 = frame (4k)
frame_vm_group_bin_18778 = frame (4k)
frame_vm_group_bin_18779 = frame (4k)
frame_vm_group_bin_1878 = frame (4k)
frame_vm_group_bin_18780 = frame (4k)
frame_vm_group_bin_18781 = frame (4k)
frame_vm_group_bin_18782 = frame (4k)
frame_vm_group_bin_18783 = frame (4k)
frame_vm_group_bin_18784 = frame (4k)
frame_vm_group_bin_18785 = frame (4k)
frame_vm_group_bin_18786 = frame (4k)
frame_vm_group_bin_18787 = frame (4k)
frame_vm_group_bin_18788 = frame (4k)
frame_vm_group_bin_18789 = frame (4k)
frame_vm_group_bin_1879 = frame (4k)
frame_vm_group_bin_18790 = frame (4k)
frame_vm_group_bin_18791 = frame (4k)
frame_vm_group_bin_18792 = frame (4k)
frame_vm_group_bin_18793 = frame (4k)
frame_vm_group_bin_18794 = frame (4k)
frame_vm_group_bin_18795 = frame (4k)
frame_vm_group_bin_18796 = frame (4k)
frame_vm_group_bin_18797 = frame (4k)
frame_vm_group_bin_18798 = frame (4k)
frame_vm_group_bin_18799 = frame (4k)
frame_vm_group_bin_1880 = frame (4k)
frame_vm_group_bin_18800 = frame (4k)
frame_vm_group_bin_18801 = frame (4k)
frame_vm_group_bin_18802 = frame (4k)
frame_vm_group_bin_18803 = frame (4k)
frame_vm_group_bin_18804 = frame (4k)
frame_vm_group_bin_18805 = frame (4k)
frame_vm_group_bin_18806 = frame (4k)
frame_vm_group_bin_18807 = frame (4k)
frame_vm_group_bin_18808 = frame (4k)
frame_vm_group_bin_18809 = frame (4k)
frame_vm_group_bin_1881 = frame (4k)
frame_vm_group_bin_18810 = frame (4k)
frame_vm_group_bin_18811 = frame (4k)
frame_vm_group_bin_18812 = frame (4k)
frame_vm_group_bin_18813 = frame (4k)
frame_vm_group_bin_18814 = frame (4k)
frame_vm_group_bin_18815 = frame (4k)
frame_vm_group_bin_18816 = frame (4k)
frame_vm_group_bin_18817 = frame (4k)
frame_vm_group_bin_18818 = frame (4k)
frame_vm_group_bin_18819 = frame (4k)
frame_vm_group_bin_1882 = frame (4k)
frame_vm_group_bin_18820 = frame (4k)
frame_vm_group_bin_18821 = frame (4k)
frame_vm_group_bin_18822 = frame (4k)
frame_vm_group_bin_18823 = frame (4k)
frame_vm_group_bin_18824 = frame (4k)
frame_vm_group_bin_18825 = frame (4k)
frame_vm_group_bin_18826 = frame (4k)
frame_vm_group_bin_18827 = frame (4k)
frame_vm_group_bin_18828 = frame (4k)
frame_vm_group_bin_18829 = frame (4k)
frame_vm_group_bin_1883 = frame (4k)
frame_vm_group_bin_18830 = frame (4k)
frame_vm_group_bin_18831 = frame (4k)
frame_vm_group_bin_18832 = frame (4k)
frame_vm_group_bin_18833 = frame (4k)
frame_vm_group_bin_18834 = frame (4k)
frame_vm_group_bin_18835 = frame (4k)
frame_vm_group_bin_18836 = frame (4k)
frame_vm_group_bin_18837 = frame (4k)
frame_vm_group_bin_18838 = frame (4k)
frame_vm_group_bin_18839 = frame (4k)
frame_vm_group_bin_1884 = frame (4k)
frame_vm_group_bin_18840 = frame (4k)
frame_vm_group_bin_18841 = frame (4k)
frame_vm_group_bin_18842 = frame (4k)
frame_vm_group_bin_18843 = frame (4k)
frame_vm_group_bin_18844 = frame (4k)
frame_vm_group_bin_18845 = frame (4k)
frame_vm_group_bin_18846 = frame (4k)
frame_vm_group_bin_18847 = frame (4k)
frame_vm_group_bin_18848 = frame (4k)
frame_vm_group_bin_18849 = frame (4k)
frame_vm_group_bin_1885 = frame (4k)
frame_vm_group_bin_18850 = frame (4k)
frame_vm_group_bin_18851 = frame (4k)
frame_vm_group_bin_18852 = frame (4k)
frame_vm_group_bin_18853 = frame (4k)
frame_vm_group_bin_18854 = frame (4k)
frame_vm_group_bin_18855 = frame (4k)
frame_vm_group_bin_18856 = frame (4k)
frame_vm_group_bin_18857 = frame (4k)
frame_vm_group_bin_18858 = frame (4k)
frame_vm_group_bin_18859 = frame (4k)
frame_vm_group_bin_1886 = frame (4k)
frame_vm_group_bin_18860 = frame (4k)
frame_vm_group_bin_18861 = frame (4k)
frame_vm_group_bin_18862 = frame (4k)
frame_vm_group_bin_18863 = frame (4k)
frame_vm_group_bin_18864 = frame (4k)
frame_vm_group_bin_18865 = frame (4k)
frame_vm_group_bin_18866 = frame (4k)
frame_vm_group_bin_18867 = frame (4k)
frame_vm_group_bin_18868 = frame (4k)
frame_vm_group_bin_18869 = frame (4k)
frame_vm_group_bin_1887 = frame (4k)
frame_vm_group_bin_18870 = frame (4k)
frame_vm_group_bin_18871 = frame (4k)
frame_vm_group_bin_18872 = frame (4k)
frame_vm_group_bin_18873 = frame (4k)
frame_vm_group_bin_18874 = frame (4k)
frame_vm_group_bin_18875 = frame (4k)
frame_vm_group_bin_18876 = frame (4k)
frame_vm_group_bin_18877 = frame (4k)
frame_vm_group_bin_18878 = frame (4k)
frame_vm_group_bin_18879 = frame (4k)
frame_vm_group_bin_1888 = frame (4k)
frame_vm_group_bin_18880 = frame (4k)
frame_vm_group_bin_18881 = frame (4k)
frame_vm_group_bin_18882 = frame (4k)
frame_vm_group_bin_18883 = frame (4k)
frame_vm_group_bin_18884 = frame (4k)
frame_vm_group_bin_18885 = frame (4k)
frame_vm_group_bin_18886 = frame (4k)
frame_vm_group_bin_18887 = frame (4k)
frame_vm_group_bin_18888 = frame (4k)
frame_vm_group_bin_18889 = frame (4k)
frame_vm_group_bin_1889 = frame (4k)
frame_vm_group_bin_18890 = frame (4k)
frame_vm_group_bin_18891 = frame (4k)
frame_vm_group_bin_18892 = frame (4k)
frame_vm_group_bin_18893 = frame (4k)
frame_vm_group_bin_18894 = frame (4k)
frame_vm_group_bin_18895 = frame (4k)
frame_vm_group_bin_18896 = frame (4k)
frame_vm_group_bin_18897 = frame (4k)
frame_vm_group_bin_18898 = frame (4k)
frame_vm_group_bin_18899 = frame (4k)
frame_vm_group_bin_1890 = frame (4k)
frame_vm_group_bin_18900 = frame (4k)
frame_vm_group_bin_18901 = frame (4k)
frame_vm_group_bin_18902 = frame (4k)
frame_vm_group_bin_18903 = frame (4k)
frame_vm_group_bin_18904 = frame (4k)
frame_vm_group_bin_18905 = frame (4k)
frame_vm_group_bin_18906 = frame (4k)
frame_vm_group_bin_18907 = frame (4k)
frame_vm_group_bin_18908 = frame (4k)
frame_vm_group_bin_18909 = frame (4k)
frame_vm_group_bin_1891 = frame (4k)
frame_vm_group_bin_18910 = frame (4k)
frame_vm_group_bin_18911 = frame (4k)
frame_vm_group_bin_18912 = frame (4k)
frame_vm_group_bin_18913 = frame (4k)
frame_vm_group_bin_18914 = frame (4k)
frame_vm_group_bin_18915 = frame (4k)
frame_vm_group_bin_18916 = frame (4k)
frame_vm_group_bin_18917 = frame (4k)
frame_vm_group_bin_18918 = frame (4k)
frame_vm_group_bin_18919 = frame (4k)
frame_vm_group_bin_1892 = frame (4k)
frame_vm_group_bin_18920 = frame (4k)
frame_vm_group_bin_18921 = frame (4k)
frame_vm_group_bin_18922 = frame (4k)
frame_vm_group_bin_18923 = frame (4k)
frame_vm_group_bin_18924 = frame (4k)
frame_vm_group_bin_18925 = frame (4k)
frame_vm_group_bin_18926 = frame (4k)
frame_vm_group_bin_18927 = frame (4k)
frame_vm_group_bin_18928 = frame (4k)
frame_vm_group_bin_18929 = frame (4k)
frame_vm_group_bin_1893 = frame (4k)
frame_vm_group_bin_18930 = frame (4k)
frame_vm_group_bin_18931 = frame (4k)
frame_vm_group_bin_18932 = frame (4k)
frame_vm_group_bin_18933 = frame (4k)
frame_vm_group_bin_18934 = frame (4k)
frame_vm_group_bin_18935 = frame (4k)
frame_vm_group_bin_18936 = frame (4k)
frame_vm_group_bin_18937 = frame (4k)
frame_vm_group_bin_18938 = frame (4k)
frame_vm_group_bin_18939 = frame (4k)
frame_vm_group_bin_1894 = frame (4k)
frame_vm_group_bin_18940 = frame (4k)
frame_vm_group_bin_18941 = frame (4k)
frame_vm_group_bin_18942 = frame (4k)
frame_vm_group_bin_18943 = frame (4k)
frame_vm_group_bin_18944 = frame (4k)
frame_vm_group_bin_18945 = frame (4k)
frame_vm_group_bin_18946 = frame (4k)
frame_vm_group_bin_18947 = frame (4k)
frame_vm_group_bin_18948 = frame (4k)
frame_vm_group_bin_18949 = frame (4k)
frame_vm_group_bin_1895 = frame (4k)
frame_vm_group_bin_18950 = frame (4k)
frame_vm_group_bin_18951 = frame (4k)
frame_vm_group_bin_18952 = frame (4k)
frame_vm_group_bin_18953 = frame (4k)
frame_vm_group_bin_18954 = frame (4k)
frame_vm_group_bin_18955 = frame (4k)
frame_vm_group_bin_18956 = frame (4k)
frame_vm_group_bin_18957 = frame (4k)
frame_vm_group_bin_18958 = frame (4k)
frame_vm_group_bin_18959 = frame (4k)
frame_vm_group_bin_1896 = frame (4k)
frame_vm_group_bin_18960 = frame (4k)
frame_vm_group_bin_18961 = frame (4k)
frame_vm_group_bin_18962 = frame (4k)
frame_vm_group_bin_18963 = frame (4k)
frame_vm_group_bin_18964 = frame (4k)
frame_vm_group_bin_18965 = frame (4k)
frame_vm_group_bin_18966 = frame (4k)
frame_vm_group_bin_18967 = frame (4k)
frame_vm_group_bin_18968 = frame (4k)
frame_vm_group_bin_18969 = frame (4k)
frame_vm_group_bin_1897 = frame (4k)
frame_vm_group_bin_18970 = frame (4k)
frame_vm_group_bin_18971 = frame (4k)
frame_vm_group_bin_18972 = frame (4k)
frame_vm_group_bin_18973 = frame (4k)
frame_vm_group_bin_18974 = frame (4k)
frame_vm_group_bin_18975 = frame (4k)
frame_vm_group_bin_18976 = frame (4k)
frame_vm_group_bin_18977 = frame (4k)
frame_vm_group_bin_18978 = frame (4k)
frame_vm_group_bin_18979 = frame (4k)
frame_vm_group_bin_1898 = frame (4k)
frame_vm_group_bin_18980 = frame (4k)
frame_vm_group_bin_18981 = frame (4k)
frame_vm_group_bin_18982 = frame (4k)
frame_vm_group_bin_18983 = frame (4k)
frame_vm_group_bin_18984 = frame (4k)
frame_vm_group_bin_18985 = frame (4k)
frame_vm_group_bin_18986 = frame (4k)
frame_vm_group_bin_18987 = frame (4k)
frame_vm_group_bin_18988 = frame (4k)
frame_vm_group_bin_18989 = frame (4k)
frame_vm_group_bin_1899 = frame (4k)
frame_vm_group_bin_18990 = frame (4k)
frame_vm_group_bin_18991 = frame (4k)
frame_vm_group_bin_18992 = frame (4k)
frame_vm_group_bin_18993 = frame (4k)
frame_vm_group_bin_18994 = frame (4k)
frame_vm_group_bin_18995 = frame (4k)
frame_vm_group_bin_18996 = frame (4k)
frame_vm_group_bin_18997 = frame (4k)
frame_vm_group_bin_18998 = frame (4k)
frame_vm_group_bin_18999 = frame (4k)
frame_vm_group_bin_1900 = frame (4k)
frame_vm_group_bin_19000 = frame (4k)
frame_vm_group_bin_19001 = frame (4k)
frame_vm_group_bin_19002 = frame (4k)
frame_vm_group_bin_19003 = frame (4k)
frame_vm_group_bin_19004 = frame (4k)
frame_vm_group_bin_19005 = frame (4k)
frame_vm_group_bin_19006 = frame (4k)
frame_vm_group_bin_19007 = frame (4k)
frame_vm_group_bin_19008 = frame (4k)
frame_vm_group_bin_19009 = frame (4k)
frame_vm_group_bin_1901 = frame (4k)
frame_vm_group_bin_19010 = frame (4k)
frame_vm_group_bin_19011 = frame (4k)
frame_vm_group_bin_19012 = frame (4k)
frame_vm_group_bin_19013 = frame (4k)
frame_vm_group_bin_19014 = frame (4k)
frame_vm_group_bin_19015 = frame (4k)
frame_vm_group_bin_19016 = frame (4k)
frame_vm_group_bin_19017 = frame (4k)
frame_vm_group_bin_19018 = frame (4k)
frame_vm_group_bin_19019 = frame (4k)
frame_vm_group_bin_1902 = frame (4k)
frame_vm_group_bin_19020 = frame (4k)
frame_vm_group_bin_19021 = frame (4k)
frame_vm_group_bin_19022 = frame (4k)
frame_vm_group_bin_19023 = frame (4k)
frame_vm_group_bin_19024 = frame (4k)
frame_vm_group_bin_19025 = frame (4k)
frame_vm_group_bin_19026 = frame (4k)
frame_vm_group_bin_19027 = frame (4k)
frame_vm_group_bin_19028 = frame (4k)
frame_vm_group_bin_19029 = frame (4k)
frame_vm_group_bin_1903 = frame (4k)
frame_vm_group_bin_19030 = frame (4k)
frame_vm_group_bin_19031 = frame (4k)
frame_vm_group_bin_19032 = frame (4k)
frame_vm_group_bin_19033 = frame (4k)
frame_vm_group_bin_19034 = frame (4k)
frame_vm_group_bin_19035 = frame (4k)
frame_vm_group_bin_19036 = frame (4k)
frame_vm_group_bin_19037 = frame (4k)
frame_vm_group_bin_19038 = frame (4k)
frame_vm_group_bin_19039 = frame (4k)
frame_vm_group_bin_1904 = frame (4k)
frame_vm_group_bin_19040 = frame (4k)
frame_vm_group_bin_19041 = frame (4k)
frame_vm_group_bin_19042 = frame (4k)
frame_vm_group_bin_19043 = frame (4k)
frame_vm_group_bin_19044 = frame (4k)
frame_vm_group_bin_19045 = frame (4k)
frame_vm_group_bin_19046 = frame (4k)
frame_vm_group_bin_19047 = frame (4k)
frame_vm_group_bin_19048 = frame (4k)
frame_vm_group_bin_19049 = frame (4k)
frame_vm_group_bin_1905 = frame (4k)
frame_vm_group_bin_19050 = frame (4k)
frame_vm_group_bin_19051 = frame (4k)
frame_vm_group_bin_19052 = frame (4k)
frame_vm_group_bin_19053 = frame (4k)
frame_vm_group_bin_19054 = frame (4k)
frame_vm_group_bin_19055 = frame (4k)
frame_vm_group_bin_19056 = frame (4k)
frame_vm_group_bin_19057 = frame (4k)
frame_vm_group_bin_19058 = frame (4k)
frame_vm_group_bin_19059 = frame (4k)
frame_vm_group_bin_1906 = frame (4k)
frame_vm_group_bin_19060 = frame (4k)
frame_vm_group_bin_19061 = frame (4k)
frame_vm_group_bin_19062 = frame (4k)
frame_vm_group_bin_19063 = frame (4k)
frame_vm_group_bin_19064 = frame (4k)
frame_vm_group_bin_19065 = frame (4k)
frame_vm_group_bin_19066 = frame (4k)
frame_vm_group_bin_19067 = frame (4k)
frame_vm_group_bin_19068 = frame (4k)
frame_vm_group_bin_19069 = frame (4k)
frame_vm_group_bin_1907 = frame (4k)
frame_vm_group_bin_19070 = frame (4k)
frame_vm_group_bin_19071 = frame (4k)
frame_vm_group_bin_19072 = frame (4k)
frame_vm_group_bin_19073 = frame (4k)
frame_vm_group_bin_19074 = frame (4k)
frame_vm_group_bin_19075 = frame (4k)
frame_vm_group_bin_19076 = frame (4k)
frame_vm_group_bin_19077 = frame (4k)
frame_vm_group_bin_19078 = frame (4k)
frame_vm_group_bin_19079 = frame (4k)
frame_vm_group_bin_1908 = frame (4k)
frame_vm_group_bin_19080 = frame (4k)
frame_vm_group_bin_19081 = frame (4k)
frame_vm_group_bin_19082 = frame (4k)
frame_vm_group_bin_19083 = frame (4k)
frame_vm_group_bin_19084 = frame (4k)
frame_vm_group_bin_19085 = frame (4k)
frame_vm_group_bin_19086 = frame (4k)
frame_vm_group_bin_19087 = frame (4k)
frame_vm_group_bin_19088 = frame (4k)
frame_vm_group_bin_19089 = frame (4k)
frame_vm_group_bin_1909 = frame (4k)
frame_vm_group_bin_19090 = frame (4k)
frame_vm_group_bin_19091 = frame (4k)
frame_vm_group_bin_19092 = frame (4k)
frame_vm_group_bin_19093 = frame (4k)
frame_vm_group_bin_19094 = frame (4k)
frame_vm_group_bin_19095 = frame (4k)
frame_vm_group_bin_19096 = frame (4k)
frame_vm_group_bin_19097 = frame (4k)
frame_vm_group_bin_19098 = frame (4k)
frame_vm_group_bin_19099 = frame (4k)
frame_vm_group_bin_1910 = frame (4k)
frame_vm_group_bin_19100 = frame (4k)
frame_vm_group_bin_19101 = frame (4k)
frame_vm_group_bin_19102 = frame (4k)
frame_vm_group_bin_19103 = frame (4k)
frame_vm_group_bin_19104 = frame (4k)
frame_vm_group_bin_19105 = frame (4k)
frame_vm_group_bin_19106 = frame (4k)
frame_vm_group_bin_19107 = frame (4k)
frame_vm_group_bin_19108 = frame (4k)
frame_vm_group_bin_19109 = frame (4k)
frame_vm_group_bin_1911 = frame (4k)
frame_vm_group_bin_19110 = frame (4k)
frame_vm_group_bin_19111 = frame (4k)
frame_vm_group_bin_19112 = frame (4k)
frame_vm_group_bin_19113 = frame (4k)
frame_vm_group_bin_19114 = frame (4k)
frame_vm_group_bin_19115 = frame (4k)
frame_vm_group_bin_19116 = frame (4k)
frame_vm_group_bin_19117 = frame (4k)
frame_vm_group_bin_19118 = frame (4k)
frame_vm_group_bin_19119 = frame (4k)
frame_vm_group_bin_1912 = frame (4k)
frame_vm_group_bin_19120 = frame (4k)
frame_vm_group_bin_19121 = frame (4k)
frame_vm_group_bin_19122 = frame (4k)
frame_vm_group_bin_19123 = frame (4k)
frame_vm_group_bin_19124 = frame (4k)
frame_vm_group_bin_19125 = frame (4k)
frame_vm_group_bin_19126 = frame (4k)
frame_vm_group_bin_19127 = frame (4k)
frame_vm_group_bin_19128 = frame (4k)
frame_vm_group_bin_19129 = frame (4k)
frame_vm_group_bin_1913 = frame (4k)
frame_vm_group_bin_19130 = frame (4k)
frame_vm_group_bin_19131 = frame (4k)
frame_vm_group_bin_19132 = frame (4k)
frame_vm_group_bin_19133 = frame (4k)
frame_vm_group_bin_19134 = frame (4k)
frame_vm_group_bin_19135 = frame (4k)
frame_vm_group_bin_19136 = frame (4k)
frame_vm_group_bin_19137 = frame (4k)
frame_vm_group_bin_19138 = frame (4k)
frame_vm_group_bin_19139 = frame (4k)
frame_vm_group_bin_1914 = frame (4k)
frame_vm_group_bin_19140 = frame (4k)
frame_vm_group_bin_19141 = frame (4k)
frame_vm_group_bin_19142 = frame (4k)
frame_vm_group_bin_19143 = frame (4k)
frame_vm_group_bin_19144 = frame (4k)
frame_vm_group_bin_19145 = frame (4k)
frame_vm_group_bin_19146 = frame (4k)
frame_vm_group_bin_19147 = frame (4k)
frame_vm_group_bin_19148 = frame (4k)
frame_vm_group_bin_19149 = frame (4k)
frame_vm_group_bin_1915 = frame (4k)
frame_vm_group_bin_19150 = frame (4k)
frame_vm_group_bin_19151 = frame (4k)
frame_vm_group_bin_19152 = frame (4k)
frame_vm_group_bin_19153 = frame (4k)
frame_vm_group_bin_19154 = frame (4k)
frame_vm_group_bin_19155 = frame (4k)
frame_vm_group_bin_19156 = frame (4k)
frame_vm_group_bin_19157 = frame (4k)
frame_vm_group_bin_19158 = frame (4k)
frame_vm_group_bin_19159 = frame (4k)
frame_vm_group_bin_1916 = frame (4k)
frame_vm_group_bin_19160 = frame (4k)
frame_vm_group_bin_19161 = frame (4k)
frame_vm_group_bin_19162 = frame (4k)
frame_vm_group_bin_19163 = frame (4k)
frame_vm_group_bin_19164 = frame (4k)
frame_vm_group_bin_19165 = frame (4k)
frame_vm_group_bin_19166 = frame (4k)
frame_vm_group_bin_19167 = frame (4k)
frame_vm_group_bin_19168 = frame (4k)
frame_vm_group_bin_19169 = frame (4k)
frame_vm_group_bin_1917 = frame (4k)
frame_vm_group_bin_19170 = frame (4k)
frame_vm_group_bin_19171 = frame (4k)
frame_vm_group_bin_19172 = frame (4k)
frame_vm_group_bin_19173 = frame (4k)
frame_vm_group_bin_19174 = frame (4k)
frame_vm_group_bin_19175 = frame (4k)
frame_vm_group_bin_19176 = frame (4k)
frame_vm_group_bin_19177 = frame (4k)
frame_vm_group_bin_19178 = frame (4k)
frame_vm_group_bin_19179 = frame (4k)
frame_vm_group_bin_1918 = frame (4k)
frame_vm_group_bin_19180 = frame (4k)
frame_vm_group_bin_19181 = frame (4k)
frame_vm_group_bin_19182 = frame (4k)
frame_vm_group_bin_19183 = frame (4k)
frame_vm_group_bin_19184 = frame (4k)
frame_vm_group_bin_19185 = frame (4k)
frame_vm_group_bin_19186 = frame (4k)
frame_vm_group_bin_19187 = frame (4k)
frame_vm_group_bin_19188 = frame (4k)
frame_vm_group_bin_19189 = frame (4k)
frame_vm_group_bin_1919 = frame (4k)
frame_vm_group_bin_19190 = frame (4k)
frame_vm_group_bin_19191 = frame (4k)
frame_vm_group_bin_19192 = frame (4k)
frame_vm_group_bin_19193 = frame (4k)
frame_vm_group_bin_19194 = frame (4k)
frame_vm_group_bin_19195 = frame (4k)
frame_vm_group_bin_19196 = frame (4k)
frame_vm_group_bin_19197 = frame (4k)
frame_vm_group_bin_19198 = frame (4k)
frame_vm_group_bin_19199 = frame (4k)
frame_vm_group_bin_1920 = frame (4k)
frame_vm_group_bin_19200 = frame (4k)
frame_vm_group_bin_19201 = frame (4k)
frame_vm_group_bin_19202 = frame (4k)
frame_vm_group_bin_19203 = frame (4k)
frame_vm_group_bin_19204 = frame (4k)
frame_vm_group_bin_19205 = frame (4k)
frame_vm_group_bin_19206 = frame (4k)
frame_vm_group_bin_19207 = frame (4k)
frame_vm_group_bin_19208 = frame (4k)
frame_vm_group_bin_19209 = frame (4k)
frame_vm_group_bin_1921 = frame (4k)
frame_vm_group_bin_19210 = frame (4k)
frame_vm_group_bin_19211 = frame (4k)
frame_vm_group_bin_19212 = frame (4k)
frame_vm_group_bin_19213 = frame (4k)
frame_vm_group_bin_19214 = frame (4k)
frame_vm_group_bin_19215 = frame (4k)
frame_vm_group_bin_19216 = frame (4k)
frame_vm_group_bin_19217 = frame (4k)
frame_vm_group_bin_19218 = frame (4k)
frame_vm_group_bin_19219 = frame (4k)
frame_vm_group_bin_1922 = frame (4k)
frame_vm_group_bin_19220 = frame (4k)
frame_vm_group_bin_19221 = frame (4k)
frame_vm_group_bin_19222 = frame (4k)
frame_vm_group_bin_19223 = frame (4k)
frame_vm_group_bin_19224 = frame (4k)
frame_vm_group_bin_19225 = frame (4k)
frame_vm_group_bin_19226 = frame (4k)
frame_vm_group_bin_19227 = frame (4k)
frame_vm_group_bin_19228 = frame (4k)
frame_vm_group_bin_19229 = frame (4k)
frame_vm_group_bin_1923 = frame (4k)
frame_vm_group_bin_19230 = frame (4k)
frame_vm_group_bin_19231 = frame (4k)
frame_vm_group_bin_19232 = frame (4k)
frame_vm_group_bin_19233 = frame (4k)
frame_vm_group_bin_19234 = frame (4k)
frame_vm_group_bin_19235 = frame (4k)
frame_vm_group_bin_19236 = frame (4k)
frame_vm_group_bin_19237 = frame (4k)
frame_vm_group_bin_19238 = frame (4k)
frame_vm_group_bin_19239 = frame (4k)
frame_vm_group_bin_1924 = frame (4k)
frame_vm_group_bin_19240 = frame (4k)
frame_vm_group_bin_19241 = frame (4k)
frame_vm_group_bin_19242 = frame (4k)
frame_vm_group_bin_19243 = frame (4k)
frame_vm_group_bin_19244 = frame (4k)
frame_vm_group_bin_19245 = frame (4k)
frame_vm_group_bin_19246 = frame (4k)
frame_vm_group_bin_19247 = frame (4k)
frame_vm_group_bin_19248 = frame (4k)
frame_vm_group_bin_19249 = frame (4k)
frame_vm_group_bin_1925 = frame (4k)
frame_vm_group_bin_19250 = frame (4k)
frame_vm_group_bin_19251 = frame (4k)
frame_vm_group_bin_19252 = frame (4k)
frame_vm_group_bin_19253 = frame (4k)
frame_vm_group_bin_19254 = frame (4k)
frame_vm_group_bin_19255 = frame (4k)
frame_vm_group_bin_19256 = frame (4k)
frame_vm_group_bin_19257 = frame (4k)
frame_vm_group_bin_19258 = frame (4k)
frame_vm_group_bin_19259 = frame (4k)
frame_vm_group_bin_1926 = frame (4k)
frame_vm_group_bin_19260 = frame (4k)
frame_vm_group_bin_19261 = frame (4k)
frame_vm_group_bin_19262 = frame (4k)
frame_vm_group_bin_19263 = frame (4k)
frame_vm_group_bin_19264 = frame (4k)
frame_vm_group_bin_19265 = frame (4k)
frame_vm_group_bin_19266 = frame (4k)
frame_vm_group_bin_19267 = frame (4k)
frame_vm_group_bin_19268 = frame (4k)
frame_vm_group_bin_19269 = frame (4k)
frame_vm_group_bin_1927 = frame (4k)
frame_vm_group_bin_19270 = frame (4k)
frame_vm_group_bin_19271 = frame (4k)
frame_vm_group_bin_19272 = frame (4k)
frame_vm_group_bin_19273 = frame (4k)
frame_vm_group_bin_19274 = frame (4k)
frame_vm_group_bin_19275 = frame (4k)
frame_vm_group_bin_19276 = frame (4k)
frame_vm_group_bin_19277 = frame (4k)
frame_vm_group_bin_19278 = frame (4k)
frame_vm_group_bin_19279 = frame (4k)
frame_vm_group_bin_1928 = frame (4k)
frame_vm_group_bin_19280 = frame (4k)
frame_vm_group_bin_19281 = frame (4k)
frame_vm_group_bin_19282 = frame (4k)
frame_vm_group_bin_19283 = frame (4k)
frame_vm_group_bin_19284 = frame (4k)
frame_vm_group_bin_19285 = frame (4k)
frame_vm_group_bin_19286 = frame (4k)
frame_vm_group_bin_19287 = frame (4k)
frame_vm_group_bin_19288 = frame (4k)
frame_vm_group_bin_19289 = frame (4k)
frame_vm_group_bin_1929 = frame (4k)
frame_vm_group_bin_19290 = frame (4k)
frame_vm_group_bin_19291 = frame (4k)
frame_vm_group_bin_19292 = frame (4k)
frame_vm_group_bin_19293 = frame (4k)
frame_vm_group_bin_19294 = frame (4k)
frame_vm_group_bin_19295 = frame (4k)
frame_vm_group_bin_19296 = frame (4k)
frame_vm_group_bin_19297 = frame (4k)
frame_vm_group_bin_19298 = frame (4k)
frame_vm_group_bin_19299 = frame (4k)
frame_vm_group_bin_1930 = frame (4k)
frame_vm_group_bin_19300 = frame (4k)
frame_vm_group_bin_19301 = frame (4k)
frame_vm_group_bin_19302 = frame (4k)
frame_vm_group_bin_19303 = frame (4k)
frame_vm_group_bin_19304 = frame (4k)
frame_vm_group_bin_19305 = frame (4k)
frame_vm_group_bin_19306 = frame (4k)
frame_vm_group_bin_19307 = frame (4k)
frame_vm_group_bin_19308 = frame (4k)
frame_vm_group_bin_19309 = frame (4k)
frame_vm_group_bin_1931 = frame (4k)
frame_vm_group_bin_19310 = frame (4k)
frame_vm_group_bin_19311 = frame (4k)
frame_vm_group_bin_19312 = frame (4k)
frame_vm_group_bin_19313 = frame (4k)
frame_vm_group_bin_19314 = frame (4k)
frame_vm_group_bin_19315 = frame (4k)
frame_vm_group_bin_19316 = frame (4k)
frame_vm_group_bin_19317 = frame (4k)
frame_vm_group_bin_19318 = frame (4k)
frame_vm_group_bin_19319 = frame (4k)
frame_vm_group_bin_1932 = frame (4k)
frame_vm_group_bin_19320 = frame (4k)
frame_vm_group_bin_19321 = frame (4k)
frame_vm_group_bin_19322 = frame (4k)
frame_vm_group_bin_19323 = frame (4k)
frame_vm_group_bin_19324 = frame (4k)
frame_vm_group_bin_19325 = frame (4k)
frame_vm_group_bin_19326 = frame (4k)
frame_vm_group_bin_19327 = frame (4k)
frame_vm_group_bin_19328 = frame (4k)
frame_vm_group_bin_19329 = frame (4k)
frame_vm_group_bin_1933 = frame (4k)
frame_vm_group_bin_19330 = frame (4k)
frame_vm_group_bin_19331 = frame (4k)
frame_vm_group_bin_19332 = frame (4k)
frame_vm_group_bin_19333 = frame (4k)
frame_vm_group_bin_19334 = frame (4k)
frame_vm_group_bin_19335 = frame (4k)
frame_vm_group_bin_19336 = frame (4k)
frame_vm_group_bin_19337 = frame (4k)
frame_vm_group_bin_19338 = frame (4k)
frame_vm_group_bin_19339 = frame (4k)
frame_vm_group_bin_1934 = frame (4k)
frame_vm_group_bin_19340 = frame (4k)
frame_vm_group_bin_19341 = frame (4k)
frame_vm_group_bin_19342 = frame (4k)
frame_vm_group_bin_19343 = frame (4k)
frame_vm_group_bin_19344 = frame (4k)
frame_vm_group_bin_19345 = frame (4k)
frame_vm_group_bin_19346 = frame (4k)
frame_vm_group_bin_19347 = frame (4k)
frame_vm_group_bin_19348 = frame (4k)
frame_vm_group_bin_19349 = frame (4k)
frame_vm_group_bin_1935 = frame (4k)
frame_vm_group_bin_19350 = frame (4k)
frame_vm_group_bin_19351 = frame (4k)
frame_vm_group_bin_19352 = frame (4k)
frame_vm_group_bin_19353 = frame (4k)
frame_vm_group_bin_19354 = frame (4k)
frame_vm_group_bin_19355 = frame (4k)
frame_vm_group_bin_19356 = frame (4k)
frame_vm_group_bin_19357 = frame (4k)
frame_vm_group_bin_19358 = frame (4k)
frame_vm_group_bin_19359 = frame (4k)
frame_vm_group_bin_1936 = frame (4k)
frame_vm_group_bin_19360 = frame (4k)
frame_vm_group_bin_19361 = frame (4k)
frame_vm_group_bin_19362 = frame (4k)
frame_vm_group_bin_19363 = frame (4k)
frame_vm_group_bin_19364 = frame (4k)
frame_vm_group_bin_19365 = frame (4k)
frame_vm_group_bin_19366 = frame (4k)
frame_vm_group_bin_19367 = frame (4k)
frame_vm_group_bin_19368 = frame (4k)
frame_vm_group_bin_19369 = frame (4k)
frame_vm_group_bin_1937 = frame (4k)
frame_vm_group_bin_19370 = frame (4k)
frame_vm_group_bin_19371 = frame (4k)
frame_vm_group_bin_19372 = frame (4k)
frame_vm_group_bin_19373 = frame (4k)
frame_vm_group_bin_19374 = frame (4k)
frame_vm_group_bin_19375 = frame (4k)
frame_vm_group_bin_19376 = frame (4k)
frame_vm_group_bin_19377 = frame (4k)
frame_vm_group_bin_19378 = frame (4k)
frame_vm_group_bin_19379 = frame (4k)
frame_vm_group_bin_1938 = frame (4k)
frame_vm_group_bin_19380 = frame (4k)
frame_vm_group_bin_19381 = frame (4k)
frame_vm_group_bin_19382 = frame (4k)
frame_vm_group_bin_19383 = frame (4k)
frame_vm_group_bin_19384 = frame (4k)
frame_vm_group_bin_19385 = frame (4k)
frame_vm_group_bin_19386 = frame (4k)
frame_vm_group_bin_19387 = frame (4k)
frame_vm_group_bin_19388 = frame (4k)
frame_vm_group_bin_19389 = frame (4k)
frame_vm_group_bin_1939 = frame (4k)
frame_vm_group_bin_19390 = frame (4k)
frame_vm_group_bin_19391 = frame (4k)
frame_vm_group_bin_19392 = frame (4k)
frame_vm_group_bin_19393 = frame (4k)
frame_vm_group_bin_19394 = frame (4k)
frame_vm_group_bin_19395 = frame (4k)
frame_vm_group_bin_19396 = frame (4k)
frame_vm_group_bin_19397 = frame (4k)
frame_vm_group_bin_19398 = frame (4k)
frame_vm_group_bin_19399 = frame (4k)
frame_vm_group_bin_1940 = frame (4k)
frame_vm_group_bin_19400 = frame (4k)
frame_vm_group_bin_19401 = frame (4k)
frame_vm_group_bin_19402 = frame (4k)
frame_vm_group_bin_19403 = frame (4k)
frame_vm_group_bin_19404 = frame (4k)
frame_vm_group_bin_19405 = frame (4k)
frame_vm_group_bin_19406 = frame (4k)
frame_vm_group_bin_19407 = frame (4k)
frame_vm_group_bin_19408 = frame (4k)
frame_vm_group_bin_19409 = frame (4k)
frame_vm_group_bin_1941 = frame (4k)
frame_vm_group_bin_19410 = frame (4k)
frame_vm_group_bin_19411 = frame (4k)
frame_vm_group_bin_19412 = frame (4k)
frame_vm_group_bin_19413 = frame (4k)
frame_vm_group_bin_19414 = frame (4k)
frame_vm_group_bin_19415 = frame (4k)
frame_vm_group_bin_19416 = frame (4k)
frame_vm_group_bin_19417 = frame (4k)
frame_vm_group_bin_19418 = frame (4k)
frame_vm_group_bin_19419 = frame (4k)
frame_vm_group_bin_1942 = frame (4k)
frame_vm_group_bin_19420 = frame (4k)
frame_vm_group_bin_19421 = frame (4k)
frame_vm_group_bin_19422 = frame (4k)
frame_vm_group_bin_19423 = frame (4k)
frame_vm_group_bin_19424 = frame (4k)
frame_vm_group_bin_19425 = frame (4k)
frame_vm_group_bin_19426 = frame (4k)
frame_vm_group_bin_19427 = frame (4k)
frame_vm_group_bin_19428 = frame (4k)
frame_vm_group_bin_19429 = frame (4k)
frame_vm_group_bin_1943 = frame (4k)
frame_vm_group_bin_19430 = frame (4k)
frame_vm_group_bin_19431 = frame (4k)
frame_vm_group_bin_19432 = frame (4k)
frame_vm_group_bin_19433 = frame (4k)
frame_vm_group_bin_19434 = frame (4k)
frame_vm_group_bin_19435 = frame (4k)
frame_vm_group_bin_19436 = frame (4k)
frame_vm_group_bin_19437 = frame (4k)
frame_vm_group_bin_19438 = frame (4k)
frame_vm_group_bin_19439 = frame (4k)
frame_vm_group_bin_1944 = frame (4k)
frame_vm_group_bin_19440 = frame (4k)
frame_vm_group_bin_19441 = frame (4k)
frame_vm_group_bin_19442 = frame (4k)
frame_vm_group_bin_19443 = frame (4k)
frame_vm_group_bin_19444 = frame (4k)
frame_vm_group_bin_19445 = frame (4k)
frame_vm_group_bin_19446 = frame (4k)
frame_vm_group_bin_19447 = frame (4k)
frame_vm_group_bin_19448 = frame (4k)
frame_vm_group_bin_19449 = frame (4k)
frame_vm_group_bin_1945 = frame (4k)
frame_vm_group_bin_19450 = frame (4k)
frame_vm_group_bin_19451 = frame (4k)
frame_vm_group_bin_19452 = frame (4k)
frame_vm_group_bin_19453 = frame (4k)
frame_vm_group_bin_19454 = frame (4k)
frame_vm_group_bin_19455 = frame (4k)
frame_vm_group_bin_19456 = frame (4k)
frame_vm_group_bin_19457 = frame (4k)
frame_vm_group_bin_19458 = frame (4k)
frame_vm_group_bin_19459 = frame (4k)
frame_vm_group_bin_1946 = frame (4k)
frame_vm_group_bin_19460 = frame (4k)
frame_vm_group_bin_19461 = frame (4k)
frame_vm_group_bin_19462 = frame (4k)
frame_vm_group_bin_19463 = frame (4k)
frame_vm_group_bin_19464 = frame (4k)
frame_vm_group_bin_19465 = frame (4k)
frame_vm_group_bin_19466 = frame (4k)
frame_vm_group_bin_19467 = frame (4k)
frame_vm_group_bin_19468 = frame (4k)
frame_vm_group_bin_19469 = frame (4k)
frame_vm_group_bin_1947 = frame (4k)
frame_vm_group_bin_19470 = frame (4k)
frame_vm_group_bin_19471 = frame (4k)
frame_vm_group_bin_19472 = frame (4k)
frame_vm_group_bin_19473 = frame (4k)
frame_vm_group_bin_19474 = frame (4k)
frame_vm_group_bin_19475 = frame (4k)
frame_vm_group_bin_19476 = frame (4k)
frame_vm_group_bin_19477 = frame (4k)
frame_vm_group_bin_19478 = frame (4k)
frame_vm_group_bin_19479 = frame (4k)
frame_vm_group_bin_1948 = frame (4k)
frame_vm_group_bin_19480 = frame (4k)
frame_vm_group_bin_19481 = frame (4k)
frame_vm_group_bin_19482 = frame (4k)
frame_vm_group_bin_19483 = frame (4k)
frame_vm_group_bin_19484 = frame (4k)
frame_vm_group_bin_19485 = frame (4k)
frame_vm_group_bin_19486 = frame (4k)
frame_vm_group_bin_19487 = frame (4k)
frame_vm_group_bin_19488 = frame (4k)
frame_vm_group_bin_19489 = frame (4k)
frame_vm_group_bin_1949 = frame (4k)
frame_vm_group_bin_19490 = frame (4k)
frame_vm_group_bin_19491 = frame (4k)
frame_vm_group_bin_19492 = frame (4k)
frame_vm_group_bin_19493 = frame (4k)
frame_vm_group_bin_19494 = frame (4k)
frame_vm_group_bin_19495 = frame (4k)
frame_vm_group_bin_19496 = frame (4k)
frame_vm_group_bin_19497 = frame (4k)
frame_vm_group_bin_19498 = frame (4k)
frame_vm_group_bin_19499 = frame (4k)
frame_vm_group_bin_1950 = frame (4k)
frame_vm_group_bin_19500 = frame (4k)
frame_vm_group_bin_19501 = frame (4k)
frame_vm_group_bin_19502 = frame (4k)
frame_vm_group_bin_19503 = frame (4k)
frame_vm_group_bin_19504 = frame (4k)
frame_vm_group_bin_19505 = frame (4k)
frame_vm_group_bin_19506 = frame (4k)
frame_vm_group_bin_19507 = frame (4k)
frame_vm_group_bin_19508 = frame (4k)
frame_vm_group_bin_19509 = frame (4k)
frame_vm_group_bin_1951 = frame (4k)
frame_vm_group_bin_19510 = frame (4k)
frame_vm_group_bin_19511 = frame (4k)
frame_vm_group_bin_19512 = frame (4k)
frame_vm_group_bin_19513 = frame (4k)
frame_vm_group_bin_19514 = frame (4k)
frame_vm_group_bin_19515 = frame (4k)
frame_vm_group_bin_19516 = frame (4k)
frame_vm_group_bin_19517 = frame (4k)
frame_vm_group_bin_19518 = frame (4k)
frame_vm_group_bin_19519 = frame (4k)
frame_vm_group_bin_1952 = frame (4k)
frame_vm_group_bin_19520 = frame (4k)
frame_vm_group_bin_19521 = frame (4k)
frame_vm_group_bin_19522 = frame (4k)
frame_vm_group_bin_19523 = frame (4k)
frame_vm_group_bin_19524 = frame (4k)
frame_vm_group_bin_19525 = frame (4k)
frame_vm_group_bin_19526 = frame (4k)
frame_vm_group_bin_19527 = frame (4k)
frame_vm_group_bin_19528 = frame (4k)
frame_vm_group_bin_19529 = frame (4k)
frame_vm_group_bin_1953 = frame (4k)
frame_vm_group_bin_19530 = frame (4k)
frame_vm_group_bin_19531 = frame (4k)
frame_vm_group_bin_19532 = frame (4k)
frame_vm_group_bin_19533 = frame (4k)
frame_vm_group_bin_19534 = frame (4k)
frame_vm_group_bin_19535 = frame (4k)
frame_vm_group_bin_19536 = frame (4k)
frame_vm_group_bin_19537 = frame (4k)
frame_vm_group_bin_19538 = frame (4k)
frame_vm_group_bin_19539 = frame (4k)
frame_vm_group_bin_1954 = frame (4k)
frame_vm_group_bin_19540 = frame (4k)
frame_vm_group_bin_19541 = frame (4k)
frame_vm_group_bin_19542 = frame (4k)
frame_vm_group_bin_19543 = frame (4k)
frame_vm_group_bin_19544 = frame (4k)
frame_vm_group_bin_19545 = frame (4k)
frame_vm_group_bin_19546 = frame (4k)
frame_vm_group_bin_19547 = frame (4k)
frame_vm_group_bin_19548 = frame (4k)
frame_vm_group_bin_19549 = frame (4k)
frame_vm_group_bin_1955 = frame (4k)
frame_vm_group_bin_19550 = frame (4k)
frame_vm_group_bin_19551 = frame (4k)
frame_vm_group_bin_19552 = frame (4k)
frame_vm_group_bin_19553 = frame (4k)
frame_vm_group_bin_19554 = frame (4k)
frame_vm_group_bin_19555 = frame (4k)
frame_vm_group_bin_19556 = frame (4k)
frame_vm_group_bin_19557 = frame (4k)
frame_vm_group_bin_19558 = frame (4k)
frame_vm_group_bin_19559 = frame (4k)
frame_vm_group_bin_1956 = frame (4k)
frame_vm_group_bin_19560 = frame (4k)
frame_vm_group_bin_19561 = frame (4k)
frame_vm_group_bin_19562 = frame (4k)
frame_vm_group_bin_19563 = frame (4k)
frame_vm_group_bin_19564 = frame (4k)
frame_vm_group_bin_19565 = frame (4k)
frame_vm_group_bin_19566 = frame (4k)
frame_vm_group_bin_19567 = frame (4k)
frame_vm_group_bin_19568 = frame (4k)
frame_vm_group_bin_19569 = frame (4k)
frame_vm_group_bin_1957 = frame (4k)
frame_vm_group_bin_19570 = frame (4k)
frame_vm_group_bin_19571 = frame (4k)
frame_vm_group_bin_19572 = frame (4k)
frame_vm_group_bin_19573 = frame (4k)
frame_vm_group_bin_19574 = frame (4k)
frame_vm_group_bin_19575 = frame (4k)
frame_vm_group_bin_19576 = frame (4k)
frame_vm_group_bin_19577 = frame (4k)
frame_vm_group_bin_19578 = frame (4k)
frame_vm_group_bin_19579 = frame (4k)
frame_vm_group_bin_1958 = frame (4k)
frame_vm_group_bin_19580 = frame (4k)
frame_vm_group_bin_19581 = frame (4k)
frame_vm_group_bin_19582 = frame (4k)
frame_vm_group_bin_19583 = frame (4k)
frame_vm_group_bin_19584 = frame (4k)
frame_vm_group_bin_19585 = frame (4k)
frame_vm_group_bin_19586 = frame (4k)
frame_vm_group_bin_19587 = frame (4k)
frame_vm_group_bin_19588 = frame (4k)
frame_vm_group_bin_19589 = frame (4k)
frame_vm_group_bin_1959 = frame (4k)
frame_vm_group_bin_19590 = frame (4k)
frame_vm_group_bin_19591 = frame (4k)
frame_vm_group_bin_19592 = frame (4k)
frame_vm_group_bin_19593 = frame (4k)
frame_vm_group_bin_19594 = frame (4k)
frame_vm_group_bin_19595 = frame (4k)
frame_vm_group_bin_19596 = frame (4k)
frame_vm_group_bin_19597 = frame (4k)
frame_vm_group_bin_19598 = frame (4k)
frame_vm_group_bin_19599 = frame (4k)
frame_vm_group_bin_1960 = frame (4k)
frame_vm_group_bin_19600 = frame (4k)
frame_vm_group_bin_19601 = frame (4k)
frame_vm_group_bin_19602 = frame (4k)
frame_vm_group_bin_19603 = frame (4k)
frame_vm_group_bin_19604 = frame (4k)
frame_vm_group_bin_19605 = frame (4k)
frame_vm_group_bin_19606 = frame (4k)
frame_vm_group_bin_19607 = frame (4k)
frame_vm_group_bin_19608 = frame (4k)
frame_vm_group_bin_19609 = frame (4k)
frame_vm_group_bin_1961 = frame (4k)
frame_vm_group_bin_19610 = frame (4k)
frame_vm_group_bin_19611 = frame (4k)
frame_vm_group_bin_19612 = frame (4k)
frame_vm_group_bin_19613 = frame (4k)
frame_vm_group_bin_19614 = frame (4k)
frame_vm_group_bin_19615 = frame (4k)
frame_vm_group_bin_19616 = frame (4k)
frame_vm_group_bin_19617 = frame (4k)
frame_vm_group_bin_19618 = frame (4k)
frame_vm_group_bin_19619 = frame (4k)
frame_vm_group_bin_1962 = frame (4k)
frame_vm_group_bin_19620 = frame (4k)
frame_vm_group_bin_19621 = frame (4k)
frame_vm_group_bin_19622 = frame (4k)
frame_vm_group_bin_19623 = frame (4k)
frame_vm_group_bin_19624 = frame (4k)
frame_vm_group_bin_19625 = frame (4k)
frame_vm_group_bin_19626 = frame (4k)
frame_vm_group_bin_19627 = frame (4k)
frame_vm_group_bin_19628 = frame (4k)
frame_vm_group_bin_19629 = frame (4k)
frame_vm_group_bin_1963 = frame (4k)
frame_vm_group_bin_19630 = frame (4k)
frame_vm_group_bin_19631 = frame (4k)
frame_vm_group_bin_19632 = frame (4k)
frame_vm_group_bin_19633 = frame (4k)
frame_vm_group_bin_19634 = frame (4k)
frame_vm_group_bin_19635 = frame (4k)
frame_vm_group_bin_19636 = frame (4k)
frame_vm_group_bin_19637 = frame (4k)
frame_vm_group_bin_19638 = frame (4k)
frame_vm_group_bin_19639 = frame (4k)
frame_vm_group_bin_1964 = frame (4k)
frame_vm_group_bin_19640 = frame (4k)
frame_vm_group_bin_19641 = frame (4k)
frame_vm_group_bin_19642 = frame (4k)
frame_vm_group_bin_19643 = frame (4k)
frame_vm_group_bin_19644 = frame (4k)
frame_vm_group_bin_19645 = frame (4k)
frame_vm_group_bin_19646 = frame (4k)
frame_vm_group_bin_19647 = frame (4k)
frame_vm_group_bin_19648 = frame (4k)
frame_vm_group_bin_19649 = frame (4k)
frame_vm_group_bin_1965 = frame (4k)
frame_vm_group_bin_19650 = frame (4k)
frame_vm_group_bin_19651 = frame (4k)
frame_vm_group_bin_19652 = frame (4k)
frame_vm_group_bin_19653 = frame (4k)
frame_vm_group_bin_19654 = frame (4k)
frame_vm_group_bin_19655 = frame (4k)
frame_vm_group_bin_19656 = frame (4k)
frame_vm_group_bin_19657 = frame (4k)
frame_vm_group_bin_19658 = frame (4k)
frame_vm_group_bin_19659 = frame (4k)
frame_vm_group_bin_1966 = frame (4k)
frame_vm_group_bin_19660 = frame (4k)
frame_vm_group_bin_19661 = frame (4k)
frame_vm_group_bin_19662 = frame (4k)
frame_vm_group_bin_19663 = frame (4k)
frame_vm_group_bin_19664 = frame (4k)
frame_vm_group_bin_19665 = frame (4k)
frame_vm_group_bin_19666 = frame (4k)
frame_vm_group_bin_19667 = frame (4k)
frame_vm_group_bin_19668 = frame (4k)
frame_vm_group_bin_19669 = frame (4k)
frame_vm_group_bin_1967 = frame (4k)
frame_vm_group_bin_19670 = frame (4k)
frame_vm_group_bin_19671 = frame (4k)
frame_vm_group_bin_19672 = frame (4k)
frame_vm_group_bin_19673 = frame (4k)
frame_vm_group_bin_19674 = frame (4k)
frame_vm_group_bin_19675 = frame (4k)
frame_vm_group_bin_19676 = frame (4k)
frame_vm_group_bin_19677 = frame (4k)
frame_vm_group_bin_19678 = frame (4k)
frame_vm_group_bin_19679 = frame (4k)
frame_vm_group_bin_1968 = frame (4k)
frame_vm_group_bin_19680 = frame (4k)
frame_vm_group_bin_19681 = frame (4k)
frame_vm_group_bin_19682 = frame (4k)
frame_vm_group_bin_19683 = frame (4k)
frame_vm_group_bin_19684 = frame (4k)
frame_vm_group_bin_19685 = frame (4k)
frame_vm_group_bin_19686 = frame (4k)
frame_vm_group_bin_19687 = frame (4k)
frame_vm_group_bin_19688 = frame (4k)
frame_vm_group_bin_19689 = frame (4k)
frame_vm_group_bin_1969 = frame (4k)
frame_vm_group_bin_19690 = frame (4k)
frame_vm_group_bin_19691 = frame (4k)
frame_vm_group_bin_19692 = frame (4k)
frame_vm_group_bin_19693 = frame (4k)
frame_vm_group_bin_19694 = frame (4k)
frame_vm_group_bin_19695 = frame (4k)
frame_vm_group_bin_19696 = frame (4k)
frame_vm_group_bin_19697 = frame (4k)
frame_vm_group_bin_19698 = frame (4k)
frame_vm_group_bin_19699 = frame (4k)
frame_vm_group_bin_1970 = frame (4k)
frame_vm_group_bin_19700 = frame (4k)
frame_vm_group_bin_19701 = frame (4k)
frame_vm_group_bin_19702 = frame (4k)
frame_vm_group_bin_19703 = frame (4k)
frame_vm_group_bin_19704 = frame (4k)
frame_vm_group_bin_19705 = frame (4k)
frame_vm_group_bin_19706 = frame (4k)
frame_vm_group_bin_19707 = frame (4k)
frame_vm_group_bin_19708 = frame (4k)
frame_vm_group_bin_19709 = frame (4k)
frame_vm_group_bin_1971 = frame (4k)
frame_vm_group_bin_19710 = frame (4k)
frame_vm_group_bin_19711 = frame (4k)
frame_vm_group_bin_19712 = frame (4k)
frame_vm_group_bin_19713 = frame (4k)
frame_vm_group_bin_19714 = frame (4k)
frame_vm_group_bin_19715 = frame (4k)
frame_vm_group_bin_19716 = frame (4k)
frame_vm_group_bin_19717 = frame (4k)
frame_vm_group_bin_19718 = frame (4k)
frame_vm_group_bin_19719 = frame (4k)
frame_vm_group_bin_1972 = frame (4k)
frame_vm_group_bin_19720 = frame (4k)
frame_vm_group_bin_19721 = frame (4k)
frame_vm_group_bin_19722 = frame (4k)
frame_vm_group_bin_19723 = frame (4k)
frame_vm_group_bin_19724 = frame (4k)
frame_vm_group_bin_19725 = frame (4k)
frame_vm_group_bin_19726 = frame (4k)
frame_vm_group_bin_19727 = frame (4k)
frame_vm_group_bin_19728 = frame (4k)
frame_vm_group_bin_19729 = frame (4k)
frame_vm_group_bin_1973 = frame (4k)
frame_vm_group_bin_19730 = frame (4k)
frame_vm_group_bin_19731 = frame (4k)
frame_vm_group_bin_19732 = frame (4k)
frame_vm_group_bin_19733 = frame (4k)
frame_vm_group_bin_19734 = frame (4k)
frame_vm_group_bin_19735 = frame (4k)
frame_vm_group_bin_19736 = frame (4k)
frame_vm_group_bin_19737 = frame (4k)
frame_vm_group_bin_19738 = frame (4k)
frame_vm_group_bin_19739 = frame (4k)
frame_vm_group_bin_1974 = frame (4k)
frame_vm_group_bin_19740 = frame (4k)
frame_vm_group_bin_19741 = frame (4k)
frame_vm_group_bin_19742 = frame (4k)
frame_vm_group_bin_19743 = frame (4k)
frame_vm_group_bin_19744 = frame (4k)
frame_vm_group_bin_19745 = frame (4k)
frame_vm_group_bin_19746 = frame (4k)
frame_vm_group_bin_19747 = frame (4k)
frame_vm_group_bin_19748 = frame (4k)
frame_vm_group_bin_19749 = frame (4k)
frame_vm_group_bin_1975 = frame (4k)
frame_vm_group_bin_19750 = frame (4k)
frame_vm_group_bin_19751 = frame (4k)
frame_vm_group_bin_19752 = frame (4k)
frame_vm_group_bin_19753 = frame (4k)
frame_vm_group_bin_19754 = frame (4k)
frame_vm_group_bin_19755 = frame (4k)
frame_vm_group_bin_19756 = frame (4k)
frame_vm_group_bin_19757 = frame (4k)
frame_vm_group_bin_19758 = frame (4k)
frame_vm_group_bin_19759 = frame (4k)
frame_vm_group_bin_1976 = frame (4k)
frame_vm_group_bin_19760 = frame (4k)
frame_vm_group_bin_19761 = frame (4k)
frame_vm_group_bin_19762 = frame (4k)
frame_vm_group_bin_19763 = frame (4k)
frame_vm_group_bin_19764 = frame (4k)
frame_vm_group_bin_19765 = frame (4k)
frame_vm_group_bin_19766 = frame (4k)
frame_vm_group_bin_19767 = frame (4k)
frame_vm_group_bin_19768 = frame (4k)
frame_vm_group_bin_19769 = frame (4k)
frame_vm_group_bin_1977 = frame (4k)
frame_vm_group_bin_19770 = frame (4k)
frame_vm_group_bin_19771 = frame (4k)
frame_vm_group_bin_19772 = frame (4k)
frame_vm_group_bin_19773 = frame (4k)
frame_vm_group_bin_19774 = frame (4k)
frame_vm_group_bin_19775 = frame (4k)
frame_vm_group_bin_19776 = frame (4k)
frame_vm_group_bin_19777 = frame (4k)
frame_vm_group_bin_19778 = frame (4k)
frame_vm_group_bin_19779 = frame (4k)
frame_vm_group_bin_1978 = frame (4k)
frame_vm_group_bin_19780 = frame (4k)
frame_vm_group_bin_19781 = frame (4k)
frame_vm_group_bin_19782 = frame (4k)
frame_vm_group_bin_19783 = frame (4k)
frame_vm_group_bin_19784 = frame (4k)
frame_vm_group_bin_19785 = frame (4k)
frame_vm_group_bin_19786 = frame (4k)
frame_vm_group_bin_19787 = frame (4k)
frame_vm_group_bin_19788 = frame (4k)
frame_vm_group_bin_19789 = frame (4k)
frame_vm_group_bin_1979 = frame (4k)
frame_vm_group_bin_19790 = frame (4k)
frame_vm_group_bin_19791 = frame (4k)
frame_vm_group_bin_19792 = frame (4k)
frame_vm_group_bin_19793 = frame (4k)
frame_vm_group_bin_19794 = frame (4k)
frame_vm_group_bin_19795 = frame (4k)
frame_vm_group_bin_19796 = frame (4k)
frame_vm_group_bin_19797 = frame (4k)
frame_vm_group_bin_19798 = frame (4k)
frame_vm_group_bin_19799 = frame (4k)
frame_vm_group_bin_1980 = frame (4k)
frame_vm_group_bin_19800 = frame (4k)
frame_vm_group_bin_19801 = frame (4k)
frame_vm_group_bin_19802 = frame (4k)
frame_vm_group_bin_19803 = frame (4k)
frame_vm_group_bin_19804 = frame (4k)
frame_vm_group_bin_19805 = frame (4k)
frame_vm_group_bin_19806 = frame (4k)
frame_vm_group_bin_19807 = frame (4k)
frame_vm_group_bin_19808 = frame (4k)
frame_vm_group_bin_19809 = frame (4k)
frame_vm_group_bin_1981 = frame (4k)
frame_vm_group_bin_19810 = frame (4k)
frame_vm_group_bin_19811 = frame (4k)
frame_vm_group_bin_19812 = frame (4k)
frame_vm_group_bin_19813 = frame (4k)
frame_vm_group_bin_19814 = frame (4k)
frame_vm_group_bin_19815 = frame (4k)
frame_vm_group_bin_19816 = frame (4k)
frame_vm_group_bin_19817 = frame (4k)
frame_vm_group_bin_19818 = frame (4k)
frame_vm_group_bin_19819 = frame (4k)
frame_vm_group_bin_1982 = frame (4k)
frame_vm_group_bin_19820 = frame (4k)
frame_vm_group_bin_19821 = frame (4k)
frame_vm_group_bin_19822 = frame (4k)
frame_vm_group_bin_19823 = frame (4k)
frame_vm_group_bin_19824 = frame (4k)
frame_vm_group_bin_19825 = frame (4k)
frame_vm_group_bin_19826 = frame (4k)
frame_vm_group_bin_19827 = frame (4k)
frame_vm_group_bin_19828 = frame (4k)
frame_vm_group_bin_19829 = frame (4k)
frame_vm_group_bin_1983 = frame (4k)
frame_vm_group_bin_19830 = frame (4k)
frame_vm_group_bin_19831 = frame (4k)
frame_vm_group_bin_19832 = frame (4k)
frame_vm_group_bin_19833 = frame (4k)
frame_vm_group_bin_19834 = frame (4k)
frame_vm_group_bin_19835 = frame (4k)
frame_vm_group_bin_19836 = frame (4k)
frame_vm_group_bin_19837 = frame (4k)
frame_vm_group_bin_19838 = frame (4k)
frame_vm_group_bin_19839 = frame (4k)
frame_vm_group_bin_1984 = frame (4k)
frame_vm_group_bin_19840 = frame (4k)
frame_vm_group_bin_19841 = frame (4k)
frame_vm_group_bin_19842 = frame (4k)
frame_vm_group_bin_19843 = frame (4k)
frame_vm_group_bin_19844 = frame (4k)
frame_vm_group_bin_19845 = frame (4k)
frame_vm_group_bin_19846 = frame (4k)
frame_vm_group_bin_19847 = frame (4k)
frame_vm_group_bin_19848 = frame (4k)
frame_vm_group_bin_19849 = frame (4k)
frame_vm_group_bin_1985 = frame (4k)
frame_vm_group_bin_19850 = frame (4k)
frame_vm_group_bin_19851 = frame (4k)
frame_vm_group_bin_19852 = frame (4k)
frame_vm_group_bin_19853 = frame (4k)
frame_vm_group_bin_19854 = frame (4k)
frame_vm_group_bin_19855 = frame (4k)
frame_vm_group_bin_19856 = frame (4k)
frame_vm_group_bin_19857 = frame (4k)
frame_vm_group_bin_19858 = frame (4k)
frame_vm_group_bin_19859 = frame (4k)
frame_vm_group_bin_1986 = frame (4k)
frame_vm_group_bin_19860 = frame (4k)
frame_vm_group_bin_19861 = frame (4k)
frame_vm_group_bin_19862 = frame (4k)
frame_vm_group_bin_19863 = frame (4k)
frame_vm_group_bin_19864 = frame (4k)
frame_vm_group_bin_19865 = frame (4k)
frame_vm_group_bin_19866 = frame (4k)
frame_vm_group_bin_19867 = frame (4k)
frame_vm_group_bin_19868 = frame (4k)
frame_vm_group_bin_19869 = frame (4k)
frame_vm_group_bin_1987 = frame (4k)
frame_vm_group_bin_19870 = frame (4k)
frame_vm_group_bin_19871 = frame (4k)
frame_vm_group_bin_19872 = frame (4k)
frame_vm_group_bin_19873 = frame (4k)
frame_vm_group_bin_19874 = frame (4k)
frame_vm_group_bin_19875 = frame (4k)
frame_vm_group_bin_19876 = frame (4k)
frame_vm_group_bin_19877 = frame (4k)
frame_vm_group_bin_19878 = frame (4k)
frame_vm_group_bin_19879 = frame (4k)
frame_vm_group_bin_1988 = frame (4k)
frame_vm_group_bin_19880 = frame (4k)
frame_vm_group_bin_19881 = frame (4k)
frame_vm_group_bin_19882 = frame (4k)
frame_vm_group_bin_19883 = frame (4k)
frame_vm_group_bin_19884 = frame (4k)
frame_vm_group_bin_19885 = frame (4k)
frame_vm_group_bin_19886 = frame (4k)
frame_vm_group_bin_19887 = frame (4k)
frame_vm_group_bin_19888 = frame (4k)
frame_vm_group_bin_19889 = frame (4k)
frame_vm_group_bin_1989 = frame (4k)
frame_vm_group_bin_19890 = frame (4k)
frame_vm_group_bin_19891 = frame (4k)
frame_vm_group_bin_19892 = frame (4k)
frame_vm_group_bin_19893 = frame (4k)
frame_vm_group_bin_19894 = frame (4k)
frame_vm_group_bin_19895 = frame (4k)
frame_vm_group_bin_19896 = frame (4k)
frame_vm_group_bin_19897 = frame (4k)
frame_vm_group_bin_19898 = frame (4k)
frame_vm_group_bin_19899 = frame (4k)
frame_vm_group_bin_1990 = frame (4k)
frame_vm_group_bin_19900 = frame (4k)
frame_vm_group_bin_19901 = frame (4k)
frame_vm_group_bin_19902 = frame (4k)
frame_vm_group_bin_19903 = frame (4k)
frame_vm_group_bin_19904 = frame (4k)
frame_vm_group_bin_19905 = frame (4k)
frame_vm_group_bin_19906 = frame (4k)
frame_vm_group_bin_19907 = frame (4k)
frame_vm_group_bin_19908 = frame (4k)
frame_vm_group_bin_19909 = frame (4k)
frame_vm_group_bin_1991 = frame (4k)
frame_vm_group_bin_19910 = frame (4k)
frame_vm_group_bin_19911 = frame (4k)
frame_vm_group_bin_19912 = frame (4k)
frame_vm_group_bin_19913 = frame (4k)
frame_vm_group_bin_19914 = frame (4k)
frame_vm_group_bin_19915 = frame (4k)
frame_vm_group_bin_19916 = frame (4k)
frame_vm_group_bin_19917 = frame (4k)
frame_vm_group_bin_19918 = frame (4k)
frame_vm_group_bin_19919 = frame (4k)
frame_vm_group_bin_1992 = frame (4k)
frame_vm_group_bin_19920 = frame (4k)
frame_vm_group_bin_19921 = frame (4k)
frame_vm_group_bin_19922 = frame (4k)
frame_vm_group_bin_19923 = frame (4k)
frame_vm_group_bin_19924 = frame (4k)
frame_vm_group_bin_19925 = frame (4k)
frame_vm_group_bin_19926 = frame (4k)
frame_vm_group_bin_19927 = frame (4k)
frame_vm_group_bin_19928 = frame (4k)
frame_vm_group_bin_19929 = frame (4k)
frame_vm_group_bin_1993 = frame (4k)
frame_vm_group_bin_19930 = frame (4k)
frame_vm_group_bin_19931 = frame (4k)
frame_vm_group_bin_19932 = frame (4k)
frame_vm_group_bin_19933 = frame (4k)
frame_vm_group_bin_19934 = frame (4k)
frame_vm_group_bin_19935 = frame (4k)
frame_vm_group_bin_19936 = frame (4k)
frame_vm_group_bin_19937 = frame (4k)
frame_vm_group_bin_19938 = frame (4k)
frame_vm_group_bin_19939 = frame (4k)
frame_vm_group_bin_1994 = frame (4k)
frame_vm_group_bin_19940 = frame (4k)
frame_vm_group_bin_19941 = frame (4k)
frame_vm_group_bin_19942 = frame (4k)
frame_vm_group_bin_19943 = frame (4k)
frame_vm_group_bin_19944 = frame (4k)
frame_vm_group_bin_19945 = frame (4k)
frame_vm_group_bin_19946 = frame (4k)
frame_vm_group_bin_19947 = frame (4k)
frame_vm_group_bin_19948 = frame (4k)
frame_vm_group_bin_19949 = frame (4k)
frame_vm_group_bin_1995 = frame (4k)
frame_vm_group_bin_19950 = frame (4k)
frame_vm_group_bin_19951 = frame (4k)
frame_vm_group_bin_19952 = frame (4k)
frame_vm_group_bin_19953 = frame (4k)
frame_vm_group_bin_19954 = frame (4k)
frame_vm_group_bin_19955 = frame (4k)
frame_vm_group_bin_19956 = frame (4k)
frame_vm_group_bin_19957 = frame (4k)
frame_vm_group_bin_19958 = frame (4k)
frame_vm_group_bin_19959 = frame (4k)
frame_vm_group_bin_1996 = frame (4k)
frame_vm_group_bin_19960 = frame (4k)
frame_vm_group_bin_19961 = frame (4k)
frame_vm_group_bin_19962 = frame (4k)
frame_vm_group_bin_19963 = frame (4k)
frame_vm_group_bin_19964 = frame (4k)
frame_vm_group_bin_19965 = frame (4k)
frame_vm_group_bin_19966 = frame (4k)
frame_vm_group_bin_19967 = frame (4k)
frame_vm_group_bin_19968 = frame (4k)
frame_vm_group_bin_19969 = frame (4k)
frame_vm_group_bin_1997 = frame (4k)
frame_vm_group_bin_19970 = frame (4k)
frame_vm_group_bin_19971 = frame (4k)
frame_vm_group_bin_19972 = frame (4k)
frame_vm_group_bin_19973 = frame (4k)
frame_vm_group_bin_19974 = frame (4k)
frame_vm_group_bin_19975 = frame (4k)
frame_vm_group_bin_19976 = frame (4k)
frame_vm_group_bin_19977 = frame (4k)
frame_vm_group_bin_19978 = frame (4k)
frame_vm_group_bin_19979 = frame (4k)
frame_vm_group_bin_1998 = frame (4k)
frame_vm_group_bin_19980 = frame (4k)
frame_vm_group_bin_19981 = frame (4k)
frame_vm_group_bin_19982 = frame (4k)
frame_vm_group_bin_19983 = frame (4k)
frame_vm_group_bin_19984 = frame (4k)
frame_vm_group_bin_19985 = frame (4k)
frame_vm_group_bin_19986 = frame (4k)
frame_vm_group_bin_19987 = frame (4k)
frame_vm_group_bin_19988 = frame (4k)
frame_vm_group_bin_19989 = frame (4k)
frame_vm_group_bin_1999 = frame (4k)
frame_vm_group_bin_19990 = frame (4k)
frame_vm_group_bin_19991 = frame (4k)
frame_vm_group_bin_19992 = frame (4k)
frame_vm_group_bin_19993 = frame (4k)
frame_vm_group_bin_19994 = frame (4k)
frame_vm_group_bin_19995 = frame (4k)
frame_vm_group_bin_19996 = frame (4k)
frame_vm_group_bin_19997 = frame (4k)
frame_vm_group_bin_19998 = frame (4k)
frame_vm_group_bin_19999 = frame (4k)
frame_vm_group_bin_2000 = frame (4k)
frame_vm_group_bin_20000 = frame (4k)
frame_vm_group_bin_20001 = frame (4k)
frame_vm_group_bin_20002 = frame (4k)
frame_vm_group_bin_20003 = frame (4k)
frame_vm_group_bin_20004 = frame (4k)
frame_vm_group_bin_20005 = frame (4k)
frame_vm_group_bin_20006 = frame (4k)
frame_vm_group_bin_20007 = frame (4k)
frame_vm_group_bin_20008 = frame (4k)
frame_vm_group_bin_20009 = frame (4k)
frame_vm_group_bin_2001 = frame (4k)
frame_vm_group_bin_20010 = frame (4k)
frame_vm_group_bin_20011 = frame (4k)
frame_vm_group_bin_20012 = frame (4k)
frame_vm_group_bin_20013 = frame (4k)
frame_vm_group_bin_20014 = frame (4k)
frame_vm_group_bin_20015 = frame (4k)
frame_vm_group_bin_20016 = frame (4k)
frame_vm_group_bin_20017 = frame (4k)
frame_vm_group_bin_20018 = frame (4k)
frame_vm_group_bin_20019 = frame (4k)
frame_vm_group_bin_2002 = frame (4k)
frame_vm_group_bin_20020 = frame (4k)
frame_vm_group_bin_20021 = frame (4k)
frame_vm_group_bin_20022 = frame (4k)
frame_vm_group_bin_20023 = frame (4k)
frame_vm_group_bin_20024 = frame (4k)
frame_vm_group_bin_20025 = frame (4k)
frame_vm_group_bin_20026 = frame (4k)
frame_vm_group_bin_20027 = frame (4k)
frame_vm_group_bin_20028 = frame (4k)
frame_vm_group_bin_20029 = frame (4k)
frame_vm_group_bin_2003 = frame (4k)
frame_vm_group_bin_20030 = frame (4k)
frame_vm_group_bin_20031 = frame (4k)
frame_vm_group_bin_20032 = frame (4k)
frame_vm_group_bin_20033 = frame (4k)
frame_vm_group_bin_20034 = frame (4k)
frame_vm_group_bin_20035 = frame (4k)
frame_vm_group_bin_20036 = frame (4k)
frame_vm_group_bin_20037 = frame (4k)
frame_vm_group_bin_20038 = frame (4k)
frame_vm_group_bin_20039 = frame (4k)
frame_vm_group_bin_2004 = frame (4k)
frame_vm_group_bin_20040 = frame (4k)
frame_vm_group_bin_20041 = frame (4k)
frame_vm_group_bin_20042 = frame (4k)
frame_vm_group_bin_20043 = frame (4k)
frame_vm_group_bin_20044 = frame (4k)
frame_vm_group_bin_20045 = frame (4k)
frame_vm_group_bin_20046 = frame (4k)
frame_vm_group_bin_20047 = frame (4k)
frame_vm_group_bin_20048 = frame (4k)
frame_vm_group_bin_20049 = frame (4k)
frame_vm_group_bin_2005 = frame (4k)
frame_vm_group_bin_20050 = frame (4k)
frame_vm_group_bin_20051 = frame (4k)
frame_vm_group_bin_20052 = frame (4k)
frame_vm_group_bin_20053 = frame (4k)
frame_vm_group_bin_20054 = frame (4k)
frame_vm_group_bin_20055 = frame (4k)
frame_vm_group_bin_20056 = frame (4k)
frame_vm_group_bin_20057 = frame (4k)
frame_vm_group_bin_20058 = frame (4k)
frame_vm_group_bin_20059 = frame (4k)
frame_vm_group_bin_2006 = frame (4k)
frame_vm_group_bin_20060 = frame (4k)
frame_vm_group_bin_20061 = frame (4k)
frame_vm_group_bin_20062 = frame (4k)
frame_vm_group_bin_20063 = frame (4k)
frame_vm_group_bin_20064 = frame (4k)
frame_vm_group_bin_20065 = frame (4k)
frame_vm_group_bin_20066 = frame (4k)
frame_vm_group_bin_20067 = frame (4k)
frame_vm_group_bin_20068 = frame (4k)
frame_vm_group_bin_20069 = frame (4k)
frame_vm_group_bin_2007 = frame (4k)
frame_vm_group_bin_20070 = frame (4k)
frame_vm_group_bin_20071 = frame (4k)
frame_vm_group_bin_20072 = frame (4k)
frame_vm_group_bin_20073 = frame (4k)
frame_vm_group_bin_20074 = frame (4k)
frame_vm_group_bin_20075 = frame (4k)
frame_vm_group_bin_20076 = frame (4k)
frame_vm_group_bin_20077 = frame (4k)
frame_vm_group_bin_20078 = frame (4k)
frame_vm_group_bin_20079 = frame (4k)
frame_vm_group_bin_2008 = frame (4k)
frame_vm_group_bin_20080 = frame (4k)
frame_vm_group_bin_20081 = frame (4k)
frame_vm_group_bin_20082 = frame (4k)
frame_vm_group_bin_20083 = frame (4k)
frame_vm_group_bin_20084 = frame (4k)
frame_vm_group_bin_20085 = frame (4k)
frame_vm_group_bin_20086 = frame (4k)
frame_vm_group_bin_20087 = frame (4k)
frame_vm_group_bin_20088 = frame (4k)
frame_vm_group_bin_20089 = frame (4k)
frame_vm_group_bin_2009 = frame (4k)
frame_vm_group_bin_20090 = frame (4k)
frame_vm_group_bin_20091 = frame (4k)
frame_vm_group_bin_20092 = frame (4k)
frame_vm_group_bin_20093 = frame (4k)
frame_vm_group_bin_20094 = frame (4k)
frame_vm_group_bin_20095 = frame (4k)
frame_vm_group_bin_20096 = frame (4k)
frame_vm_group_bin_20097 = frame (4k)
frame_vm_group_bin_20098 = frame (4k)
frame_vm_group_bin_20099 = frame (4k)
frame_vm_group_bin_2010 = frame (4k)
frame_vm_group_bin_20100 = frame (4k)
frame_vm_group_bin_20101 = frame (4k)
frame_vm_group_bin_20102 = frame (4k)
frame_vm_group_bin_20103 = frame (4k)
frame_vm_group_bin_20104 = frame (4k)
frame_vm_group_bin_20105 = frame (4k)
frame_vm_group_bin_20106 = frame (4k)
frame_vm_group_bin_20107 = frame (4k)
frame_vm_group_bin_20108 = frame (4k)
frame_vm_group_bin_20109 = frame (4k)
frame_vm_group_bin_2011 = frame (4k)
frame_vm_group_bin_20110 = frame (4k)
frame_vm_group_bin_20111 = frame (4k)
frame_vm_group_bin_20112 = frame (4k)
frame_vm_group_bin_20113 = frame (4k)
frame_vm_group_bin_20114 = frame (4k)
frame_vm_group_bin_20115 = frame (4k)
frame_vm_group_bin_20116 = frame (4k)
frame_vm_group_bin_20117 = frame (4k)
frame_vm_group_bin_20118 = frame (4k)
frame_vm_group_bin_20119 = frame (4k)
frame_vm_group_bin_2012 = frame (4k)
frame_vm_group_bin_20120 = frame (4k)
frame_vm_group_bin_20121 = frame (4k)
frame_vm_group_bin_20122 = frame (4k)
frame_vm_group_bin_20123 = frame (4k)
frame_vm_group_bin_20124 = frame (4k)
frame_vm_group_bin_20125 = frame (4k)
frame_vm_group_bin_20126 = frame (4k)
frame_vm_group_bin_20127 = frame (4k)
frame_vm_group_bin_20128 = frame (4k)
frame_vm_group_bin_20129 = frame (4k)
frame_vm_group_bin_2013 = frame (4k)
frame_vm_group_bin_20130 = frame (4k)
frame_vm_group_bin_20131 = frame (4k)
frame_vm_group_bin_20132 = frame (4k)
frame_vm_group_bin_20133 = frame (4k)
frame_vm_group_bin_20134 = frame (4k)
frame_vm_group_bin_20135 = frame (4k)
frame_vm_group_bin_20136 = frame (4k)
frame_vm_group_bin_20137 = frame (4k)
frame_vm_group_bin_20138 = frame (4k)
frame_vm_group_bin_20139 = frame (4k)
frame_vm_group_bin_2014 = frame (4k)
frame_vm_group_bin_20140 = frame (4k)
frame_vm_group_bin_20141 = frame (4k)
frame_vm_group_bin_20142 = frame (4k)
frame_vm_group_bin_20143 = frame (4k)
frame_vm_group_bin_20144 = frame (4k)
frame_vm_group_bin_20145 = frame (4k)
frame_vm_group_bin_20146 = frame (4k)
frame_vm_group_bin_20147 = frame (4k)
frame_vm_group_bin_20148 = frame (4k)
frame_vm_group_bin_20149 = frame (4k)
frame_vm_group_bin_2015 = frame (4k)
frame_vm_group_bin_20150 = frame (4k)
frame_vm_group_bin_20151 = frame (4k)
frame_vm_group_bin_20152 = frame (4k)
frame_vm_group_bin_20153 = frame (4k)
frame_vm_group_bin_20154 = frame (4k)
frame_vm_group_bin_20155 = frame (4k)
frame_vm_group_bin_20156 = frame (4k)
frame_vm_group_bin_20157 = frame (4k)
frame_vm_group_bin_20158 = frame (4k)
frame_vm_group_bin_20159 = frame (4k)
frame_vm_group_bin_2016 = frame (4k)
frame_vm_group_bin_20160 = frame (4k)
frame_vm_group_bin_20161 = frame (4k)
frame_vm_group_bin_20162 = frame (4k)
frame_vm_group_bin_20163 = frame (4k)
frame_vm_group_bin_20164 = frame (4k)
frame_vm_group_bin_20165 = frame (4k)
frame_vm_group_bin_20166 = frame (4k)
frame_vm_group_bin_20167 = frame (4k)
frame_vm_group_bin_20168 = frame (4k)
frame_vm_group_bin_20169 = frame (4k)
frame_vm_group_bin_2017 = frame (4k)
frame_vm_group_bin_20170 = frame (4k)
frame_vm_group_bin_20171 = frame (4k)
frame_vm_group_bin_20172 = frame (4k)
frame_vm_group_bin_20173 = frame (4k)
frame_vm_group_bin_20174 = frame (4k)
frame_vm_group_bin_20175 = frame (4k)
frame_vm_group_bin_20176 = frame (4k)
frame_vm_group_bin_20177 = frame (4k)
frame_vm_group_bin_20178 = frame (4k)
frame_vm_group_bin_20179 = frame (4k)
frame_vm_group_bin_2018 = frame (4k)
frame_vm_group_bin_20180 = frame (4k)
frame_vm_group_bin_20181 = frame (4k)
frame_vm_group_bin_20182 = frame (4k)
frame_vm_group_bin_20183 = frame (4k)
frame_vm_group_bin_20184 = frame (4k)
frame_vm_group_bin_20185 = frame (4k)
frame_vm_group_bin_20186 = frame (4k)
frame_vm_group_bin_20187 = frame (4k)
frame_vm_group_bin_20188 = frame (4k)
frame_vm_group_bin_20189 = frame (4k)
frame_vm_group_bin_2019 = frame (4k)
frame_vm_group_bin_20190 = frame (4k)
frame_vm_group_bin_20191 = frame (4k)
frame_vm_group_bin_20192 = frame (4k)
frame_vm_group_bin_20193 = frame (4k)
frame_vm_group_bin_20194 = frame (4k)
frame_vm_group_bin_20195 = frame (4k)
frame_vm_group_bin_20196 = frame (4k)
frame_vm_group_bin_20197 = frame (4k)
frame_vm_group_bin_20198 = frame (4k)
frame_vm_group_bin_20199 = frame (4k)
frame_vm_group_bin_2020 = frame (4k)
frame_vm_group_bin_20200 = frame (4k)
frame_vm_group_bin_20201 = frame (4k)
frame_vm_group_bin_20202 = frame (4k)
frame_vm_group_bin_20203 = frame (4k)
frame_vm_group_bin_20204 = frame (4k)
frame_vm_group_bin_20205 = frame (4k)
frame_vm_group_bin_20206 = frame (4k)
frame_vm_group_bin_20207 = frame (4k)
frame_vm_group_bin_20208 = frame (4k)
frame_vm_group_bin_20209 = frame (4k)
frame_vm_group_bin_2021 = frame (4k)
frame_vm_group_bin_20210 = frame (4k)
frame_vm_group_bin_20211 = frame (4k)
frame_vm_group_bin_20212 = frame (4k)
frame_vm_group_bin_20213 = frame (4k)
frame_vm_group_bin_20214 = frame (4k)
frame_vm_group_bin_20215 = frame (4k)
frame_vm_group_bin_20216 = frame (4k)
frame_vm_group_bin_20217 = frame (4k)
frame_vm_group_bin_20218 = frame (4k)
frame_vm_group_bin_20219 = frame (4k)
frame_vm_group_bin_2022 = frame (4k)
frame_vm_group_bin_20220 = frame (4k)
frame_vm_group_bin_20221 = frame (4k)
frame_vm_group_bin_20222 = frame (4k)
frame_vm_group_bin_20223 = frame (4k)
frame_vm_group_bin_20224 = frame (4k)
frame_vm_group_bin_20225 = frame (4k)
frame_vm_group_bin_20226 = frame (4k)
frame_vm_group_bin_20227 = frame (4k)
frame_vm_group_bin_20228 = frame (4k)
frame_vm_group_bin_20229 = frame (4k)
frame_vm_group_bin_2023 = frame (4k)
frame_vm_group_bin_20230 = frame (4k)
frame_vm_group_bin_20231 = frame (4k)
frame_vm_group_bin_20232 = frame (4k)
frame_vm_group_bin_20233 = frame (4k)
frame_vm_group_bin_20234 = frame (4k)
frame_vm_group_bin_20235 = frame (4k)
frame_vm_group_bin_20236 = frame (4k)
frame_vm_group_bin_20237 = frame (4k)
frame_vm_group_bin_20238 = frame (4k)
frame_vm_group_bin_20239 = frame (4k)
frame_vm_group_bin_2024 = frame (4k)
frame_vm_group_bin_20240 = frame (4k)
frame_vm_group_bin_20241 = frame (4k)
frame_vm_group_bin_20242 = frame (4k)
frame_vm_group_bin_20243 = frame (4k)
frame_vm_group_bin_20244 = frame (4k)
frame_vm_group_bin_20245 = frame (4k)
frame_vm_group_bin_20246 = frame (4k)
frame_vm_group_bin_20247 = frame (4k)
frame_vm_group_bin_20248 = frame (4k)
frame_vm_group_bin_20249 = frame (4k)
frame_vm_group_bin_2025 = frame (4k)
frame_vm_group_bin_20250 = frame (4k)
frame_vm_group_bin_20251 = frame (4k)
frame_vm_group_bin_20252 = frame (4k)
frame_vm_group_bin_20253 = frame (4k)
frame_vm_group_bin_20254 = frame (4k)
frame_vm_group_bin_20255 = frame (4k)
frame_vm_group_bin_20256 = frame (4k)
frame_vm_group_bin_20257 = frame (4k)
frame_vm_group_bin_20258 = frame (4k)
frame_vm_group_bin_20259 = frame (4k)
frame_vm_group_bin_2026 = frame (4k)
frame_vm_group_bin_20260 = frame (4k)
frame_vm_group_bin_20261 = frame (4k)
frame_vm_group_bin_20262 = frame (4k)
frame_vm_group_bin_20263 = frame (4k)
frame_vm_group_bin_20264 = frame (4k)
frame_vm_group_bin_20265 = frame (4k)
frame_vm_group_bin_20266 = frame (4k)
frame_vm_group_bin_20267 = frame (4k)
frame_vm_group_bin_20268 = frame (4k)
frame_vm_group_bin_20269 = frame (4k)
frame_vm_group_bin_2027 = frame (4k)
frame_vm_group_bin_20270 = frame (4k)
frame_vm_group_bin_20271 = frame (4k)
frame_vm_group_bin_20272 = frame (4k)
frame_vm_group_bin_20273 = frame (4k)
frame_vm_group_bin_20274 = frame (4k)
frame_vm_group_bin_20275 = frame (4k)
frame_vm_group_bin_20276 = frame (4k)
frame_vm_group_bin_20277 = frame (4k)
frame_vm_group_bin_20278 = frame (4k)
frame_vm_group_bin_20279 = frame (4k)
frame_vm_group_bin_2028 = frame (4k)
frame_vm_group_bin_20280 = frame (4k)
frame_vm_group_bin_20281 = frame (4k)
frame_vm_group_bin_20282 = frame (4k)
frame_vm_group_bin_20283 = frame (4k)
frame_vm_group_bin_20284 = frame (4k)
frame_vm_group_bin_20285 = frame (4k)
frame_vm_group_bin_20286 = frame (4k)
frame_vm_group_bin_20287 = frame (4k)
frame_vm_group_bin_20288 = frame (4k)
frame_vm_group_bin_20289 = frame (4k)
frame_vm_group_bin_2029 = frame (4k)
frame_vm_group_bin_20290 = frame (4k)
frame_vm_group_bin_20291 = frame (4k)
frame_vm_group_bin_20292 = frame (4k)
frame_vm_group_bin_20293 = frame (4k)
frame_vm_group_bin_20294 = frame (4k)
frame_vm_group_bin_20295 = frame (4k)
frame_vm_group_bin_20296 = frame (4k)
frame_vm_group_bin_20297 = frame (4k)
frame_vm_group_bin_20298 = frame (4k)
frame_vm_group_bin_20299 = frame (4k)
frame_vm_group_bin_2030 = frame (4k)
frame_vm_group_bin_20300 = frame (4k)
frame_vm_group_bin_20301 = frame (4k)
frame_vm_group_bin_20302 = frame (4k)
frame_vm_group_bin_20303 = frame (4k)
frame_vm_group_bin_20304 = frame (4k)
frame_vm_group_bin_20305 = frame (4k)
frame_vm_group_bin_20306 = frame (4k)
frame_vm_group_bin_20307 = frame (4k)
frame_vm_group_bin_20308 = frame (4k)
frame_vm_group_bin_20309 = frame (4k)
frame_vm_group_bin_2031 = frame (4k)
frame_vm_group_bin_20310 = frame (4k)
frame_vm_group_bin_20311 = frame (4k)
frame_vm_group_bin_20312 = frame (4k)
frame_vm_group_bin_20313 = frame (4k)
frame_vm_group_bin_20314 = frame (4k)
frame_vm_group_bin_20315 = frame (4k)
frame_vm_group_bin_20316 = frame (4k)
frame_vm_group_bin_20317 = frame (4k)
frame_vm_group_bin_20318 = frame (4k)
frame_vm_group_bin_20319 = frame (4k)
frame_vm_group_bin_2032 = frame (4k)
frame_vm_group_bin_20320 = frame (4k)
frame_vm_group_bin_20321 = frame (4k)
frame_vm_group_bin_20322 = frame (4k)
frame_vm_group_bin_20323 = frame (4k)
frame_vm_group_bin_20324 = frame (4k)
frame_vm_group_bin_20325 = frame (4k)
frame_vm_group_bin_20326 = frame (4k)
frame_vm_group_bin_20327 = frame (4k)
frame_vm_group_bin_20328 = frame (4k)
frame_vm_group_bin_20329 = frame (4k)
frame_vm_group_bin_2033 = frame (4k)
frame_vm_group_bin_20330 = frame (4k)
frame_vm_group_bin_20331 = frame (4k)
frame_vm_group_bin_20332 = frame (4k)
frame_vm_group_bin_20333 = frame (4k)
frame_vm_group_bin_20334 = frame (4k)
frame_vm_group_bin_20335 = frame (4k)
frame_vm_group_bin_20336 = frame (4k)
frame_vm_group_bin_20337 = frame (4k)
frame_vm_group_bin_20338 = frame (4k)
frame_vm_group_bin_20339 = frame (4k)
frame_vm_group_bin_2034 = frame (4k)
frame_vm_group_bin_20340 = frame (4k)
frame_vm_group_bin_20341 = frame (4k)
frame_vm_group_bin_20342 = frame (4k)
frame_vm_group_bin_20343 = frame (4k)
frame_vm_group_bin_20344 = frame (4k)
frame_vm_group_bin_20345 = frame (4k)
frame_vm_group_bin_20346 = frame (4k)
frame_vm_group_bin_20347 = frame (4k)
frame_vm_group_bin_20348 = frame (4k)
frame_vm_group_bin_20349 = frame (4k)
frame_vm_group_bin_2035 = frame (4k)
frame_vm_group_bin_20350 = frame (4k)
frame_vm_group_bin_20351 = frame (4k)
frame_vm_group_bin_20352 = frame (4k)
frame_vm_group_bin_20353 = frame (4k)
frame_vm_group_bin_20354 = frame (4k)
frame_vm_group_bin_20355 = frame (4k)
frame_vm_group_bin_20356 = frame (4k)
frame_vm_group_bin_20357 = frame (4k)
frame_vm_group_bin_20358 = frame (4k)
frame_vm_group_bin_20359 = frame (4k)
frame_vm_group_bin_2036 = frame (4k)
frame_vm_group_bin_20360 = frame (4k)
frame_vm_group_bin_20361 = frame (4k)
frame_vm_group_bin_20362 = frame (4k)
frame_vm_group_bin_20363 = frame (4k)
frame_vm_group_bin_20364 = frame (4k)
frame_vm_group_bin_20365 = frame (4k)
frame_vm_group_bin_20366 = frame (4k)
frame_vm_group_bin_20367 = frame (4k)
frame_vm_group_bin_20368 = frame (4k)
frame_vm_group_bin_20369 = frame (4k)
frame_vm_group_bin_2037 = frame (4k)
frame_vm_group_bin_20370 = frame (4k)
frame_vm_group_bin_20371 = frame (4k)
frame_vm_group_bin_20372 = frame (4k)
frame_vm_group_bin_20373 = frame (4k)
frame_vm_group_bin_20374 = frame (4k)
frame_vm_group_bin_20375 = frame (4k)
frame_vm_group_bin_20376 = frame (4k)
frame_vm_group_bin_20377 = frame (4k)
frame_vm_group_bin_20378 = frame (4k)
frame_vm_group_bin_20379 = frame (4k)
frame_vm_group_bin_2038 = frame (4k)
frame_vm_group_bin_20380 = frame (4k)
frame_vm_group_bin_20381 = frame (4k)
frame_vm_group_bin_20382 = frame (4k)
frame_vm_group_bin_20383 = frame (4k)
frame_vm_group_bin_20384 = frame (4k)
frame_vm_group_bin_20385 = frame (4k)
frame_vm_group_bin_20386 = frame (4k)
frame_vm_group_bin_20387 = frame (4k)
frame_vm_group_bin_20388 = frame (4k)
frame_vm_group_bin_20389 = frame (4k)
frame_vm_group_bin_2039 = frame (4k)
frame_vm_group_bin_20390 = frame (4k)
frame_vm_group_bin_20391 = frame (4k)
frame_vm_group_bin_20392 = frame (4k)
frame_vm_group_bin_20393 = frame (4k)
frame_vm_group_bin_20394 = frame (4k)
frame_vm_group_bin_20395 = frame (4k)
frame_vm_group_bin_20396 = frame (4k)
frame_vm_group_bin_20397 = frame (4k)
frame_vm_group_bin_20398 = frame (4k)
frame_vm_group_bin_20399 = frame (4k)
frame_vm_group_bin_2040 = frame (4k)
frame_vm_group_bin_20400 = frame (4k)
frame_vm_group_bin_20401 = frame (4k)
frame_vm_group_bin_20402 = frame (4k)
frame_vm_group_bin_20403 = frame (4k)
frame_vm_group_bin_20404 = frame (4k)
frame_vm_group_bin_20405 = frame (4k)
frame_vm_group_bin_20406 = frame (4k)
frame_vm_group_bin_20407 = frame (4k)
frame_vm_group_bin_20408 = frame (4k)
frame_vm_group_bin_20409 = frame (4k)
frame_vm_group_bin_2041 = frame (4k)
frame_vm_group_bin_20410 = frame (4k)
frame_vm_group_bin_20411 = frame (4k)
frame_vm_group_bin_20412 = frame (4k)
frame_vm_group_bin_20413 = frame (4k)
frame_vm_group_bin_20414 = frame (4k)
frame_vm_group_bin_20415 = frame (4k)
frame_vm_group_bin_20416 = frame (4k)
frame_vm_group_bin_20417 = frame (4k)
frame_vm_group_bin_20418 = frame (4k)
frame_vm_group_bin_20419 = frame (4k)
frame_vm_group_bin_2042 = frame (4k)
frame_vm_group_bin_20420 = frame (4k)
frame_vm_group_bin_20421 = frame (4k)
frame_vm_group_bin_20422 = frame (4k)
frame_vm_group_bin_20423 = frame (4k)
frame_vm_group_bin_20424 = frame (4k)
frame_vm_group_bin_20425 = frame (4k)
frame_vm_group_bin_20426 = frame (4k)
frame_vm_group_bin_20427 = frame (4k)
frame_vm_group_bin_20428 = frame (4k)
frame_vm_group_bin_20429 = frame (4k)
frame_vm_group_bin_2043 = frame (4k)
frame_vm_group_bin_20430 = frame (4k)
frame_vm_group_bin_20431 = frame (4k)
frame_vm_group_bin_20432 = frame (4k)
frame_vm_group_bin_20433 = frame (4k)
frame_vm_group_bin_20434 = frame (4k)
frame_vm_group_bin_20435 = frame (4k)
frame_vm_group_bin_20436 = frame (4k)
frame_vm_group_bin_20437 = frame (4k)
frame_vm_group_bin_20438 = frame (4k)
frame_vm_group_bin_20439 = frame (4k)
frame_vm_group_bin_2044 = frame (4k)
frame_vm_group_bin_20440 = frame (4k)
frame_vm_group_bin_20441 = frame (4k)
frame_vm_group_bin_20442 = frame (4k)
frame_vm_group_bin_20443 = frame (4k)
frame_vm_group_bin_20444 = frame (4k)
frame_vm_group_bin_20445 = frame (4k)
frame_vm_group_bin_20446 = frame (4k)
frame_vm_group_bin_20447 = frame (4k)
frame_vm_group_bin_20448 = frame (4k)
frame_vm_group_bin_20449 = frame (4k)
frame_vm_group_bin_2045 = frame (4k)
frame_vm_group_bin_20450 = frame (4k)
frame_vm_group_bin_20451 = frame (4k)
frame_vm_group_bin_20452 = frame (4k)
frame_vm_group_bin_20453 = frame (4k)
frame_vm_group_bin_20454 = frame (4k)
frame_vm_group_bin_20455 = frame (4k)
frame_vm_group_bin_20456 = frame (4k)
frame_vm_group_bin_20457 = frame (4k)
frame_vm_group_bin_20458 = frame (4k)
frame_vm_group_bin_20459 = frame (4k)
frame_vm_group_bin_2046 = frame (4k)
frame_vm_group_bin_20460 = frame (4k)
frame_vm_group_bin_20461 = frame (4k)
frame_vm_group_bin_20462 = frame (4k)
frame_vm_group_bin_20463 = frame (4k)
frame_vm_group_bin_20464 = frame (4k)
frame_vm_group_bin_20465 = frame (4k)
frame_vm_group_bin_20466 = frame (4k)
frame_vm_group_bin_20467 = frame (4k)
frame_vm_group_bin_20468 = frame (4k)
frame_vm_group_bin_20469 = frame (4k)
frame_vm_group_bin_2047 = frame (4k)
frame_vm_group_bin_20470 = frame (4k)
frame_vm_group_bin_20471 = frame (4k)
frame_vm_group_bin_20472 = frame (4k)
frame_vm_group_bin_20473 = frame (4k)
frame_vm_group_bin_20474 = frame (4k)
frame_vm_group_bin_20475 = frame (4k)
frame_vm_group_bin_20476 = frame (4k)
frame_vm_group_bin_20477 = frame (4k)
frame_vm_group_bin_20478 = frame (4k)
frame_vm_group_bin_20479 = frame (4k)
frame_vm_group_bin_2048 = frame (4k)
frame_vm_group_bin_20480 = frame (4k)
frame_vm_group_bin_20481 = frame (4k)
frame_vm_group_bin_20482 = frame (4k)
frame_vm_group_bin_20483 = frame (4k)
frame_vm_group_bin_20484 = frame (4k)
frame_vm_group_bin_20485 = frame (4k)
frame_vm_group_bin_20486 = frame (4k)
frame_vm_group_bin_20487 = frame (4k)
frame_vm_group_bin_20488 = frame (4k)
frame_vm_group_bin_20489 = frame (4k)
frame_vm_group_bin_2049 = frame (4k)
frame_vm_group_bin_20490 = frame (4k)
frame_vm_group_bin_20491 = frame (4k)
frame_vm_group_bin_20492 = frame (4k)
frame_vm_group_bin_20493 = frame (4k)
frame_vm_group_bin_20494 = frame (4k)
frame_vm_group_bin_20495 = frame (4k)
frame_vm_group_bin_20496 = frame (4k)
frame_vm_group_bin_20497 = frame (4k)
frame_vm_group_bin_20498 = frame (4k)
frame_vm_group_bin_20499 = frame (4k)
frame_vm_group_bin_2050 = frame (4k)
frame_vm_group_bin_20500 = frame (4k)
frame_vm_group_bin_20501 = frame (4k)
frame_vm_group_bin_20502 = frame (4k)
frame_vm_group_bin_20503 = frame (4k)
frame_vm_group_bin_20504 = frame (4k)
frame_vm_group_bin_20505 = frame (4k)
frame_vm_group_bin_20506 = frame (4k)
frame_vm_group_bin_20507 = frame (4k)
frame_vm_group_bin_20508 = frame (4k)
frame_vm_group_bin_20509 = frame (4k)
frame_vm_group_bin_2051 = frame (4k)
frame_vm_group_bin_20510 = frame (4k)
frame_vm_group_bin_20511 = frame (4k)
frame_vm_group_bin_20512 = frame (4k)
frame_vm_group_bin_20513 = frame (4k)
frame_vm_group_bin_20514 = frame (4k)
frame_vm_group_bin_20515 = frame (4k)
frame_vm_group_bin_20516 = frame (4k)
frame_vm_group_bin_20517 = frame (4k)
frame_vm_group_bin_20518 = frame (4k)
frame_vm_group_bin_20519 = frame (4k)
frame_vm_group_bin_2052 = frame (4k)
frame_vm_group_bin_20520 = frame (4k)
frame_vm_group_bin_20521 = frame (4k)
frame_vm_group_bin_20522 = frame (4k)
frame_vm_group_bin_20523 = frame (4k)
frame_vm_group_bin_20524 = frame (4k)
frame_vm_group_bin_20525 = frame (4k)
frame_vm_group_bin_20526 = frame (4k)
frame_vm_group_bin_20527 = frame (4k)
frame_vm_group_bin_20528 = frame (4k)
frame_vm_group_bin_20529 = frame (4k)
frame_vm_group_bin_2053 = frame (4k)
frame_vm_group_bin_20530 = frame (4k)
frame_vm_group_bin_20531 = frame (4k)
frame_vm_group_bin_20532 = frame (4k)
frame_vm_group_bin_20533 = frame (4k)
frame_vm_group_bin_20534 = frame (4k)
frame_vm_group_bin_20535 = frame (4k)
frame_vm_group_bin_20536 = frame (4k)
frame_vm_group_bin_20537 = frame (4k)
frame_vm_group_bin_20538 = frame (4k)
frame_vm_group_bin_20539 = frame (4k)
frame_vm_group_bin_2054 = frame (4k)
frame_vm_group_bin_20540 = frame (4k)
frame_vm_group_bin_20541 = frame (4k)
frame_vm_group_bin_20542 = frame (4k)
frame_vm_group_bin_20543 = frame (4k)
frame_vm_group_bin_20544 = frame (4k)
frame_vm_group_bin_20545 = frame (4k)
frame_vm_group_bin_20546 = frame (4k)
frame_vm_group_bin_20547 = frame (4k)
frame_vm_group_bin_20548 = frame (4k)
frame_vm_group_bin_20549 = frame (4k)
frame_vm_group_bin_2055 = frame (4k)
frame_vm_group_bin_20550 = frame (4k)
frame_vm_group_bin_20551 = frame (4k)
frame_vm_group_bin_20552 = frame (4k)
frame_vm_group_bin_20553 = frame (4k)
frame_vm_group_bin_20554 = frame (4k)
frame_vm_group_bin_20555 = frame (4k)
frame_vm_group_bin_20556 = frame (4k)
frame_vm_group_bin_20557 = frame (4k)
frame_vm_group_bin_20558 = frame (4k)
frame_vm_group_bin_20559 = frame (4k)
frame_vm_group_bin_2056 = frame (4k)
frame_vm_group_bin_20560 = frame (4k)
frame_vm_group_bin_20561 = frame (4k)
frame_vm_group_bin_20562 = frame (4k)
frame_vm_group_bin_20563 = frame (4k)
frame_vm_group_bin_20564 = frame (4k)
frame_vm_group_bin_20565 = frame (4k)
frame_vm_group_bin_20566 = frame (4k)
frame_vm_group_bin_20567 = frame (4k)
frame_vm_group_bin_20568 = frame (4k)
frame_vm_group_bin_20569 = frame (4k)
frame_vm_group_bin_2057 = frame (4k)
frame_vm_group_bin_20570 = frame (4k)
frame_vm_group_bin_20571 = frame (4k)
frame_vm_group_bin_20572 = frame (4k)
frame_vm_group_bin_20573 = frame (4k)
frame_vm_group_bin_20574 = frame (4k)
frame_vm_group_bin_20575 = frame (4k)
frame_vm_group_bin_20576 = frame (4k)
frame_vm_group_bin_20577 = frame (4k)
frame_vm_group_bin_20578 = frame (4k)
frame_vm_group_bin_20579 = frame (4k)
frame_vm_group_bin_2058 = frame (4k)
frame_vm_group_bin_20580 = frame (4k)
frame_vm_group_bin_20581 = frame (4k)
frame_vm_group_bin_20582 = frame (4k)
frame_vm_group_bin_20583 = frame (4k)
frame_vm_group_bin_20584 = frame (4k)
frame_vm_group_bin_20585 = frame (4k)
frame_vm_group_bin_20586 = frame (4k)
frame_vm_group_bin_20587 = frame (4k)
frame_vm_group_bin_20588 = frame (4k)
frame_vm_group_bin_20589 = frame (4k)
frame_vm_group_bin_2059 = frame (4k)
frame_vm_group_bin_20590 = frame (4k)
frame_vm_group_bin_20591 = frame (4k)
frame_vm_group_bin_20592 = frame (4k)
frame_vm_group_bin_20593 = frame (4k)
frame_vm_group_bin_20594 = frame (4k)
frame_vm_group_bin_20595 = frame (4k)
frame_vm_group_bin_20596 = frame (4k)
frame_vm_group_bin_20597 = frame (4k)
frame_vm_group_bin_20598 = frame (4k)
frame_vm_group_bin_20599 = frame (4k)
frame_vm_group_bin_2060 = frame (4k)
frame_vm_group_bin_20600 = frame (4k)
frame_vm_group_bin_20601 = frame (4k)
frame_vm_group_bin_20602 = frame (4k)
frame_vm_group_bin_20603 = frame (4k)
frame_vm_group_bin_20604 = frame (4k)
frame_vm_group_bin_20605 = frame (4k)
frame_vm_group_bin_20606 = frame (4k)
frame_vm_group_bin_20607 = frame (4k)
frame_vm_group_bin_20608 = frame (4k)
frame_vm_group_bin_20609 = frame (4k)
frame_vm_group_bin_2061 = frame (4k)
frame_vm_group_bin_20610 = frame (4k)
frame_vm_group_bin_20611 = frame (4k)
frame_vm_group_bin_20612 = frame (4k)
frame_vm_group_bin_20613 = frame (4k)
frame_vm_group_bin_20614 = frame (4k)
frame_vm_group_bin_20615 = frame (4k)
frame_vm_group_bin_20616 = frame (4k)
frame_vm_group_bin_20617 = frame (4k)
frame_vm_group_bin_20618 = frame (4k)
frame_vm_group_bin_20619 = frame (4k)
frame_vm_group_bin_2062 = frame (4k)
frame_vm_group_bin_20620 = frame (4k)
frame_vm_group_bin_20621 = frame (4k)
frame_vm_group_bin_20622 = frame (4k)
frame_vm_group_bin_20623 = frame (4k)
frame_vm_group_bin_20624 = frame (4k)
frame_vm_group_bin_20625 = frame (4k)
frame_vm_group_bin_20626 = frame (4k)
frame_vm_group_bin_20627 = frame (4k)
frame_vm_group_bin_20628 = frame (4k)
frame_vm_group_bin_20629 = frame (4k)
frame_vm_group_bin_2063 = frame (4k)
frame_vm_group_bin_20630 = frame (4k)
frame_vm_group_bin_20631 = frame (4k)
frame_vm_group_bin_20632 = frame (4k)
frame_vm_group_bin_20633 = frame (4k)
frame_vm_group_bin_20634 = frame (4k)
frame_vm_group_bin_20635 = frame (4k)
frame_vm_group_bin_20636 = frame (4k)
frame_vm_group_bin_20637 = frame (4k)
frame_vm_group_bin_20638 = frame (4k)
frame_vm_group_bin_20639 = frame (4k)
frame_vm_group_bin_2064 = frame (4k)
frame_vm_group_bin_20640 = frame (4k)
frame_vm_group_bin_20641 = frame (4k)
frame_vm_group_bin_20642 = frame (4k)
frame_vm_group_bin_20643 = frame (4k)
frame_vm_group_bin_20644 = frame (4k)
frame_vm_group_bin_20645 = frame (4k)
frame_vm_group_bin_20646 = frame (4k)
frame_vm_group_bin_20647 = frame (4k)
frame_vm_group_bin_20648 = frame (4k)
frame_vm_group_bin_20649 = frame (4k)
frame_vm_group_bin_2065 = frame (4k)
frame_vm_group_bin_20650 = frame (4k)
frame_vm_group_bin_20651 = frame (4k)
frame_vm_group_bin_20652 = frame (4k)
frame_vm_group_bin_20653 = frame (4k)
frame_vm_group_bin_20654 = frame (4k)
frame_vm_group_bin_20655 = frame (4k)
frame_vm_group_bin_20656 = frame (4k)
frame_vm_group_bin_20657 = frame (4k)
frame_vm_group_bin_20658 = frame (4k)
frame_vm_group_bin_20659 = frame (4k)
frame_vm_group_bin_2066 = frame (4k)
frame_vm_group_bin_20660 = frame (4k)
frame_vm_group_bin_20661 = frame (4k)
frame_vm_group_bin_20662 = frame (4k)
frame_vm_group_bin_20663 = frame (4k)
frame_vm_group_bin_20664 = frame (4k)
frame_vm_group_bin_20665 = frame (4k)
frame_vm_group_bin_20666 = frame (4k)
frame_vm_group_bin_20667 = frame (4k)
frame_vm_group_bin_20668 = frame (4k)
frame_vm_group_bin_20669 = frame (4k)
frame_vm_group_bin_2067 = frame (4k)
frame_vm_group_bin_20670 = frame (4k)
frame_vm_group_bin_20671 = frame (4k)
frame_vm_group_bin_20672 = frame (4k)
frame_vm_group_bin_20673 = frame (4k)
frame_vm_group_bin_20674 = frame (4k)
frame_vm_group_bin_20675 = frame (4k)
frame_vm_group_bin_20676 = frame (4k)
frame_vm_group_bin_20677 = frame (4k)
frame_vm_group_bin_20678 = frame (4k)
frame_vm_group_bin_20679 = frame (4k)
frame_vm_group_bin_2068 = frame (4k)
frame_vm_group_bin_20680 = frame (4k)
frame_vm_group_bin_20681 = frame (4k)
frame_vm_group_bin_20682 = frame (4k)
frame_vm_group_bin_20683 = frame (4k)
frame_vm_group_bin_20684 = frame (4k)
frame_vm_group_bin_20685 = frame (4k)
frame_vm_group_bin_20686 = frame (4k)
frame_vm_group_bin_20687 = frame (4k)
frame_vm_group_bin_20688 = frame (4k)
frame_vm_group_bin_20689 = frame (4k)
frame_vm_group_bin_2069 = frame (4k)
frame_vm_group_bin_20690 = frame (4k)
frame_vm_group_bin_20691 = frame (4k)
frame_vm_group_bin_20692 = frame (4k)
frame_vm_group_bin_20693 = frame (4k)
frame_vm_group_bin_20694 = frame (4k)
frame_vm_group_bin_20695 = frame (4k)
frame_vm_group_bin_20696 = frame (4k)
frame_vm_group_bin_20697 = frame (4k)
frame_vm_group_bin_20698 = frame (4k)
frame_vm_group_bin_20699 = frame (4k)
frame_vm_group_bin_2070 = frame (4k)
frame_vm_group_bin_20700 = frame (4k)
frame_vm_group_bin_20701 = frame (4k)
frame_vm_group_bin_20702 = frame (4k)
frame_vm_group_bin_20703 = frame (4k)
frame_vm_group_bin_20704 = frame (4k)
frame_vm_group_bin_20705 = frame (4k)
frame_vm_group_bin_20706 = frame (4k)
frame_vm_group_bin_20707 = frame (4k)
frame_vm_group_bin_20708 = frame (4k)
frame_vm_group_bin_20709 = frame (4k)
frame_vm_group_bin_2071 = frame (4k)
frame_vm_group_bin_20710 = frame (4k)
frame_vm_group_bin_20711 = frame (4k)
frame_vm_group_bin_20712 = frame (4k)
frame_vm_group_bin_20713 = frame (4k)
frame_vm_group_bin_20714 = frame (4k)
frame_vm_group_bin_20715 = frame (4k)
frame_vm_group_bin_20716 = frame (4k)
frame_vm_group_bin_20717 = frame (4k)
frame_vm_group_bin_20718 = frame (4k)
frame_vm_group_bin_20719 = frame (4k)
frame_vm_group_bin_2072 = frame (4k)
frame_vm_group_bin_20720 = frame (4k)
frame_vm_group_bin_20721 = frame (4k)
frame_vm_group_bin_20722 = frame (4k)
frame_vm_group_bin_20723 = frame (4k)
frame_vm_group_bin_20724 = frame (4k)
frame_vm_group_bin_20725 = frame (4k)
frame_vm_group_bin_20726 = frame (4k)
frame_vm_group_bin_20727 = frame (4k)
frame_vm_group_bin_20728 = frame (4k)
frame_vm_group_bin_20729 = frame (4k)
frame_vm_group_bin_2073 = frame (4k)
frame_vm_group_bin_20730 = frame (4k)
frame_vm_group_bin_20731 = frame (4k)
frame_vm_group_bin_20732 = frame (4k)
frame_vm_group_bin_20733 = frame (4k)
frame_vm_group_bin_20734 = frame (4k)
frame_vm_group_bin_20735 = frame (4k)
frame_vm_group_bin_20736 = frame (4k)
frame_vm_group_bin_20737 = frame (4k)
frame_vm_group_bin_20738 = frame (4k)
frame_vm_group_bin_20739 = frame (4k)
frame_vm_group_bin_2074 = frame (4k)
frame_vm_group_bin_20740 = frame (4k)
frame_vm_group_bin_20741 = frame (4k)
frame_vm_group_bin_20742 = frame (4k)
frame_vm_group_bin_20743 = frame (4k)
frame_vm_group_bin_20744 = frame (4k)
frame_vm_group_bin_20745 = frame (4k)
frame_vm_group_bin_20746 = frame (4k)
frame_vm_group_bin_20747 = frame (4k)
frame_vm_group_bin_20748 = frame (4k)
frame_vm_group_bin_20749 = frame (4k)
frame_vm_group_bin_2075 = frame (4k)
frame_vm_group_bin_20750 = frame (4k)
frame_vm_group_bin_20751 = frame (4k)
frame_vm_group_bin_20752 = frame (4k)
frame_vm_group_bin_20753 = frame (4k)
frame_vm_group_bin_20754 = frame (4k)
frame_vm_group_bin_20755 = frame (4k)
frame_vm_group_bin_20756 = frame (4k)
frame_vm_group_bin_20757 = frame (4k)
frame_vm_group_bin_20758 = frame (4k)
frame_vm_group_bin_20759 = frame (4k)
frame_vm_group_bin_2076 = frame (4k)
frame_vm_group_bin_20760 = frame (4k)
frame_vm_group_bin_20761 = frame (4k)
frame_vm_group_bin_20762 = frame (4k)
frame_vm_group_bin_20763 = frame (4k)
frame_vm_group_bin_20764 = frame (4k)
frame_vm_group_bin_20765 = frame (4k)
frame_vm_group_bin_20766 = frame (4k)
frame_vm_group_bin_20767 = frame (4k)
frame_vm_group_bin_20768 = frame (4k)
frame_vm_group_bin_20769 = frame (4k)
frame_vm_group_bin_2077 = frame (4k)
frame_vm_group_bin_20770 = frame (4k)
frame_vm_group_bin_20771 = frame (4k)
frame_vm_group_bin_20772 = frame (4k)
frame_vm_group_bin_20773 = frame (4k)
frame_vm_group_bin_20774 = frame (4k)
frame_vm_group_bin_20775 = frame (4k)
frame_vm_group_bin_20776 = frame (4k)
frame_vm_group_bin_20777 = frame (4k)
frame_vm_group_bin_20778 = frame (4k)
frame_vm_group_bin_20779 = frame (4k)
frame_vm_group_bin_2078 = frame (4k)
frame_vm_group_bin_20780 = frame (4k)
frame_vm_group_bin_20781 = frame (4k)
frame_vm_group_bin_20782 = frame (4k)
frame_vm_group_bin_20783 = frame (4k)
frame_vm_group_bin_20784 = frame (4k)
frame_vm_group_bin_20785 = frame (4k)
frame_vm_group_bin_20786 = frame (4k)
frame_vm_group_bin_20787 = frame (4k)
frame_vm_group_bin_20788 = frame (4k)
frame_vm_group_bin_20789 = frame (4k)
frame_vm_group_bin_2079 = frame (4k)
frame_vm_group_bin_20790 = frame (4k)
frame_vm_group_bin_20791 = frame (4k)
frame_vm_group_bin_20792 = frame (4k)
frame_vm_group_bin_20793 = frame (4k)
frame_vm_group_bin_20794 = frame (4k)
frame_vm_group_bin_20795 = frame (4k)
frame_vm_group_bin_20796 = frame (4k)
frame_vm_group_bin_20797 = frame (4k)
frame_vm_group_bin_20798 = frame (4k)
frame_vm_group_bin_20799 = frame (4k)
frame_vm_group_bin_2080 = frame (4k)
frame_vm_group_bin_20800 = frame (4k)
frame_vm_group_bin_20801 = frame (4k)
frame_vm_group_bin_20802 = frame (4k)
frame_vm_group_bin_20803 = frame (4k)
frame_vm_group_bin_20804 = frame (4k)
frame_vm_group_bin_20805 = frame (4k)
frame_vm_group_bin_20806 = frame (4k)
frame_vm_group_bin_20807 = frame (4k)
frame_vm_group_bin_20808 = frame (4k)
frame_vm_group_bin_20809 = frame (4k)
frame_vm_group_bin_2081 = frame (4k)
frame_vm_group_bin_20810 = frame (4k)
frame_vm_group_bin_20811 = frame (4k)
frame_vm_group_bin_20812 = frame (4k)
frame_vm_group_bin_20813 = frame (4k)
frame_vm_group_bin_20814 = frame (4k)
frame_vm_group_bin_20815 = frame (4k)
frame_vm_group_bin_20816 = frame (4k)
frame_vm_group_bin_20817 = frame (4k)
frame_vm_group_bin_20818 = frame (4k)
frame_vm_group_bin_20819 = frame (4k)
frame_vm_group_bin_2082 = frame (4k)
frame_vm_group_bin_20820 = frame (4k)
frame_vm_group_bin_20821 = frame (4k)
frame_vm_group_bin_20822 = frame (4k)
frame_vm_group_bin_20823 = frame (4k)
frame_vm_group_bin_20824 = frame (4k)
frame_vm_group_bin_20825 = frame (4k)
frame_vm_group_bin_20826 = frame (4k)
frame_vm_group_bin_20827 = frame (4k)
frame_vm_group_bin_20828 = frame (4k)
frame_vm_group_bin_20829 = frame (4k)
frame_vm_group_bin_2083 = frame (4k)
frame_vm_group_bin_20830 = frame (4k)
frame_vm_group_bin_20831 = frame (4k)
frame_vm_group_bin_20832 = frame (4k)
frame_vm_group_bin_20833 = frame (4k)
frame_vm_group_bin_20834 = frame (4k)
frame_vm_group_bin_20835 = frame (4k)
frame_vm_group_bin_20836 = frame (4k)
frame_vm_group_bin_20837 = frame (4k)
frame_vm_group_bin_20838 = frame (4k)
frame_vm_group_bin_20839 = frame (4k)
frame_vm_group_bin_2084 = frame (4k)
frame_vm_group_bin_20840 = frame (4k)
frame_vm_group_bin_20841 = frame (4k)
frame_vm_group_bin_20842 = frame (4k)
frame_vm_group_bin_20843 = frame (4k)
frame_vm_group_bin_20844 = frame (4k)
frame_vm_group_bin_20845 = frame (4k)
frame_vm_group_bin_20846 = frame (4k)
frame_vm_group_bin_20847 = frame (4k)
frame_vm_group_bin_20848 = frame (4k)
frame_vm_group_bin_20849 = frame (4k)
frame_vm_group_bin_2085 = frame (4k)
frame_vm_group_bin_20850 = frame (4k)
frame_vm_group_bin_20851 = frame (4k)
frame_vm_group_bin_20852 = frame (4k)
frame_vm_group_bin_20853 = frame (4k)
frame_vm_group_bin_20854 = frame (4k)
frame_vm_group_bin_20855 = frame (4k)
frame_vm_group_bin_20856 = frame (4k)
frame_vm_group_bin_20857 = frame (4k)
frame_vm_group_bin_20858 = frame (4k)
frame_vm_group_bin_20859 = frame (4k)
frame_vm_group_bin_2086 = frame (4k)
frame_vm_group_bin_20860 = frame (4k)
frame_vm_group_bin_20861 = frame (4k)
frame_vm_group_bin_20862 = frame (4k)
frame_vm_group_bin_20863 = frame (4k)
frame_vm_group_bin_20864 = frame (4k)
frame_vm_group_bin_20865 = frame (4k)
frame_vm_group_bin_20866 = frame (4k)
frame_vm_group_bin_20867 = frame (4k)
frame_vm_group_bin_20868 = frame (4k)
frame_vm_group_bin_20869 = frame (4k)
frame_vm_group_bin_2087 = frame (4k)
frame_vm_group_bin_20870 = frame (4k)
frame_vm_group_bin_20871 = frame (4k)
frame_vm_group_bin_20872 = frame (4k)
frame_vm_group_bin_20873 = frame (4k)
frame_vm_group_bin_20874 = frame (4k)
frame_vm_group_bin_20875 = frame (4k)
frame_vm_group_bin_20876 = frame (4k)
frame_vm_group_bin_20877 = frame (4k)
frame_vm_group_bin_20878 = frame (4k)
frame_vm_group_bin_20879 = frame (4k)
frame_vm_group_bin_2088 = frame (4k)
frame_vm_group_bin_20880 = frame (4k)
frame_vm_group_bin_20881 = frame (4k)
frame_vm_group_bin_20882 = frame (4k)
frame_vm_group_bin_20883 = frame (4k)
frame_vm_group_bin_20884 = frame (4k)
frame_vm_group_bin_20885 = frame (4k)
frame_vm_group_bin_20886 = frame (4k)
frame_vm_group_bin_20887 = frame (4k)
frame_vm_group_bin_20888 = frame (4k)
frame_vm_group_bin_20889 = frame (4k)
frame_vm_group_bin_2089 = frame (4k)
frame_vm_group_bin_20890 = frame (4k)
frame_vm_group_bin_20891 = frame (4k)
frame_vm_group_bin_20892 = frame (4k)
frame_vm_group_bin_20893 = frame (4k)
frame_vm_group_bin_20894 = frame (4k)
frame_vm_group_bin_20895 = frame (4k)
frame_vm_group_bin_20896 = frame (4k)
frame_vm_group_bin_20897 = frame (4k)
frame_vm_group_bin_20898 = frame (4k)
frame_vm_group_bin_20899 = frame (4k)
frame_vm_group_bin_2090 = frame (4k)
frame_vm_group_bin_20900 = frame (4k)
frame_vm_group_bin_20901 = frame (4k)
frame_vm_group_bin_20902 = frame (4k)
frame_vm_group_bin_20903 = frame (4k)
frame_vm_group_bin_20904 = frame (4k)
frame_vm_group_bin_20905 = frame (4k)
frame_vm_group_bin_20906 = frame (4k)
frame_vm_group_bin_20907 = frame (4k)
frame_vm_group_bin_20908 = frame (4k)
frame_vm_group_bin_20909 = frame (4k)
frame_vm_group_bin_2091 = frame (4k)
frame_vm_group_bin_20910 = frame (4k)
frame_vm_group_bin_20911 = frame (4k)
frame_vm_group_bin_20912 = frame (4k)
frame_vm_group_bin_20913 = frame (4k)
frame_vm_group_bin_20914 = frame (4k)
frame_vm_group_bin_20915 = frame (4k)
frame_vm_group_bin_20916 = frame (4k)
frame_vm_group_bin_20917 = frame (4k)
frame_vm_group_bin_20918 = frame (4k)
frame_vm_group_bin_20919 = frame (4k)
frame_vm_group_bin_2092 = frame (4k)
frame_vm_group_bin_20920 = frame (4k)
frame_vm_group_bin_20921 = frame (4k)
frame_vm_group_bin_20922 = frame (4k)
frame_vm_group_bin_20923 = frame (4k)
frame_vm_group_bin_20924 = frame (4k)
frame_vm_group_bin_20925 = frame (4k)
frame_vm_group_bin_20926 = frame (4k)
frame_vm_group_bin_20927 = frame (4k)
frame_vm_group_bin_20928 = frame (4k)
frame_vm_group_bin_20929 = frame (4k)
frame_vm_group_bin_2093 = frame (4k)
frame_vm_group_bin_20930 = frame (4k)
frame_vm_group_bin_20931 = frame (4k)
frame_vm_group_bin_20932 = frame (4k)
frame_vm_group_bin_20933 = frame (4k)
frame_vm_group_bin_20934 = frame (4k)
frame_vm_group_bin_20935 = frame (4k)
frame_vm_group_bin_20936 = frame (4k)
frame_vm_group_bin_20937 = frame (4k)
frame_vm_group_bin_20938 = frame (4k)
frame_vm_group_bin_20939 = frame (4k)
frame_vm_group_bin_2094 = frame (4k)
frame_vm_group_bin_20940 = frame (4k)
frame_vm_group_bin_20941 = frame (4k)
frame_vm_group_bin_20942 = frame (4k)
frame_vm_group_bin_20943 = frame (4k)
frame_vm_group_bin_20944 = frame (4k)
frame_vm_group_bin_20945 = frame (4k)
frame_vm_group_bin_20946 = frame (4k)
frame_vm_group_bin_20947 = frame (4k)
frame_vm_group_bin_20948 = frame (4k)
frame_vm_group_bin_20949 = frame (4k)
frame_vm_group_bin_2095 = frame (4k)
frame_vm_group_bin_20950 = frame (4k)
frame_vm_group_bin_20951 = frame (4k)
frame_vm_group_bin_20952 = frame (4k)
frame_vm_group_bin_20953 = frame (4k)
frame_vm_group_bin_20954 = frame (4k)
frame_vm_group_bin_20955 = frame (4k)
frame_vm_group_bin_20956 = frame (4k)
frame_vm_group_bin_20957 = frame (4k)
frame_vm_group_bin_20958 = frame (4k)
frame_vm_group_bin_20959 = frame (4k)
frame_vm_group_bin_2096 = frame (4k)
frame_vm_group_bin_20960 = frame (4k)
frame_vm_group_bin_20961 = frame (4k)
frame_vm_group_bin_20962 = frame (4k)
frame_vm_group_bin_20963 = frame (4k)
frame_vm_group_bin_20964 = frame (4k)
frame_vm_group_bin_20965 = frame (4k)
frame_vm_group_bin_20966 = frame (4k)
frame_vm_group_bin_20967 = frame (4k)
frame_vm_group_bin_20968 = frame (4k)
frame_vm_group_bin_20969 = frame (4k)
frame_vm_group_bin_2097 = frame (4k)
frame_vm_group_bin_20970 = frame (4k)
frame_vm_group_bin_20971 = frame (4k)
frame_vm_group_bin_20972 = frame (4k)
frame_vm_group_bin_20973 = frame (4k)
frame_vm_group_bin_20974 = frame (4k)
frame_vm_group_bin_20975 = frame (4k)
frame_vm_group_bin_20976 = frame (4k)
frame_vm_group_bin_20977 = frame (4k)
frame_vm_group_bin_20978 = frame (4k)
frame_vm_group_bin_20979 = frame (4k)
frame_vm_group_bin_2098 = frame (4k)
frame_vm_group_bin_20980 = frame (4k)
frame_vm_group_bin_20981 = frame (4k)
frame_vm_group_bin_20982 = frame (4k)
frame_vm_group_bin_20983 = frame (4k)
frame_vm_group_bin_20984 = frame (4k)
frame_vm_group_bin_20985 = frame (4k)
frame_vm_group_bin_20986 = frame (4k)
frame_vm_group_bin_20987 = frame (4k)
frame_vm_group_bin_20988 = frame (4k)
frame_vm_group_bin_20989 = frame (4k)
frame_vm_group_bin_2099 = frame (4k)
frame_vm_group_bin_20990 = frame (4k)
frame_vm_group_bin_20991 = frame (4k)
frame_vm_group_bin_20992 = frame (4k)
frame_vm_group_bin_20993 = frame (4k)
frame_vm_group_bin_20994 = frame (4k)
frame_vm_group_bin_20995 = frame (4k)
frame_vm_group_bin_20996 = frame (4k)
frame_vm_group_bin_20997 = frame (4k)
frame_vm_group_bin_20998 = frame (4k)
frame_vm_group_bin_20999 = frame (4k)
frame_vm_group_bin_2100 = frame (4k)
frame_vm_group_bin_21000 = frame (4k)
frame_vm_group_bin_21001 = frame (4k)
frame_vm_group_bin_21002 = frame (4k)
frame_vm_group_bin_21003 = frame (4k)
frame_vm_group_bin_21004 = frame (4k)
frame_vm_group_bin_21005 = frame (4k)
frame_vm_group_bin_21006 = frame (4k)
frame_vm_group_bin_21007 = frame (4k)
frame_vm_group_bin_21008 = frame (4k)
frame_vm_group_bin_21009 = frame (4k)
frame_vm_group_bin_2101 = frame (4k)
frame_vm_group_bin_21010 = frame (4k)
frame_vm_group_bin_21011 = frame (4k)
frame_vm_group_bin_21012 = frame (4k)
frame_vm_group_bin_21013 = frame (4k)
frame_vm_group_bin_21014 = frame (4k)
frame_vm_group_bin_21015 = frame (4k)
frame_vm_group_bin_21016 = frame (4k)
frame_vm_group_bin_21017 = frame (4k)
frame_vm_group_bin_21018 = frame (4k)
frame_vm_group_bin_21019 = frame (4k)
frame_vm_group_bin_2102 = frame (4k)
frame_vm_group_bin_21020 = frame (4k)
frame_vm_group_bin_21021 = frame (4k)
frame_vm_group_bin_21022 = frame (4k)
frame_vm_group_bin_21023 = frame (4k)
frame_vm_group_bin_21024 = frame (4k)
frame_vm_group_bin_21025 = frame (4k)
frame_vm_group_bin_21026 = frame (4k)
frame_vm_group_bin_21027 = frame (4k)
frame_vm_group_bin_21028 = frame (4k)
frame_vm_group_bin_21029 = frame (4k)
frame_vm_group_bin_2103 = frame (4k)
frame_vm_group_bin_21030 = frame (4k)
frame_vm_group_bin_21031 = frame (4k)
frame_vm_group_bin_21032 = frame (4k)
frame_vm_group_bin_21033 = frame (4k)
frame_vm_group_bin_21034 = frame (4k)
frame_vm_group_bin_21035 = frame (4k)
frame_vm_group_bin_21036 = frame (4k)
frame_vm_group_bin_21037 = frame (4k)
frame_vm_group_bin_21038 = frame (4k)
frame_vm_group_bin_21039 = frame (4k)
frame_vm_group_bin_2104 = frame (4k)
frame_vm_group_bin_21040 = frame (4k)
frame_vm_group_bin_21041 = frame (4k)
frame_vm_group_bin_21042 = frame (4k)
frame_vm_group_bin_21043 = frame (4k)
frame_vm_group_bin_21044 = frame (4k)
frame_vm_group_bin_21045 = frame (4k)
frame_vm_group_bin_21046 = frame (4k)
frame_vm_group_bin_21047 = frame (4k)
frame_vm_group_bin_21048 = frame (4k)
frame_vm_group_bin_21049 = frame (4k)
frame_vm_group_bin_2105 = frame (4k)
frame_vm_group_bin_21050 = frame (4k)
frame_vm_group_bin_21051 = frame (4k)
frame_vm_group_bin_21052 = frame (4k)
frame_vm_group_bin_21053 = frame (4k)
frame_vm_group_bin_21054 = frame (4k)
frame_vm_group_bin_21055 = frame (4k)
frame_vm_group_bin_21056 = frame (4k)
frame_vm_group_bin_21057 = frame (4k)
frame_vm_group_bin_21058 = frame (4k)
frame_vm_group_bin_21059 = frame (4k)
frame_vm_group_bin_2106 = frame (4k)
frame_vm_group_bin_21060 = frame (4k)
frame_vm_group_bin_21061 = frame (4k)
frame_vm_group_bin_21062 = frame (4k)
frame_vm_group_bin_21063 = frame (4k)
frame_vm_group_bin_21064 = frame (4k)
frame_vm_group_bin_21065 = frame (4k)
frame_vm_group_bin_21066 = frame (4k)
frame_vm_group_bin_21067 = frame (4k)
frame_vm_group_bin_21068 = frame (4k)
frame_vm_group_bin_21069 = frame (4k)
frame_vm_group_bin_2107 = frame (4k)
frame_vm_group_bin_21070 = frame (4k)
frame_vm_group_bin_21071 = frame (4k)
frame_vm_group_bin_21072 = frame (4k)
frame_vm_group_bin_21073 = frame (4k)
frame_vm_group_bin_21074 = frame (4k)
frame_vm_group_bin_21075 = frame (4k)
frame_vm_group_bin_21076 = frame (4k)
frame_vm_group_bin_21077 = frame (4k)
frame_vm_group_bin_21078 = frame (4k)
frame_vm_group_bin_21079 = frame (4k)
frame_vm_group_bin_2108 = frame (4k)
frame_vm_group_bin_21080 = frame (4k)
frame_vm_group_bin_21081 = frame (4k)
frame_vm_group_bin_21082 = frame (4k)
frame_vm_group_bin_21083 = frame (4k)
frame_vm_group_bin_21084 = frame (4k)
frame_vm_group_bin_21085 = frame (4k)
frame_vm_group_bin_21086 = frame (4k)
frame_vm_group_bin_21087 = frame (4k)
frame_vm_group_bin_21088 = frame (4k)
frame_vm_group_bin_21089 = frame (4k)
frame_vm_group_bin_2109 = frame (4k)
frame_vm_group_bin_21090 = frame (4k)
frame_vm_group_bin_21091 = frame (4k)
frame_vm_group_bin_21092 = frame (4k)
frame_vm_group_bin_21093 = frame (4k)
frame_vm_group_bin_21094 = frame (4k)
frame_vm_group_bin_21095 = frame (4k)
frame_vm_group_bin_21096 = frame (4k)
frame_vm_group_bin_21097 = frame (4k)
frame_vm_group_bin_21098 = frame (4k)
frame_vm_group_bin_21099 = frame (4k)
frame_vm_group_bin_2110 = frame (4k)
frame_vm_group_bin_21100 = frame (4k)
frame_vm_group_bin_21101 = frame (4k)
frame_vm_group_bin_21102 = frame (4k)
frame_vm_group_bin_21103 = frame (4k)
frame_vm_group_bin_21104 = frame (4k)
frame_vm_group_bin_21105 = frame (4k)
frame_vm_group_bin_21106 = frame (4k)
frame_vm_group_bin_21107 = frame (4k)
frame_vm_group_bin_21108 = frame (4k)
frame_vm_group_bin_21109 = frame (4k)
frame_vm_group_bin_2111 = frame (4k)
frame_vm_group_bin_21110 = frame (4k)
frame_vm_group_bin_21111 = frame (4k)
frame_vm_group_bin_21112 = frame (4k)
frame_vm_group_bin_21113 = frame (4k)
frame_vm_group_bin_21114 = frame (4k)
frame_vm_group_bin_21115 = frame (4k)
frame_vm_group_bin_21116 = frame (4k)
frame_vm_group_bin_21117 = frame (4k)
frame_vm_group_bin_21118 = frame (4k)
frame_vm_group_bin_21119 = frame (4k)
frame_vm_group_bin_2112 = frame (4k)
frame_vm_group_bin_21120 = frame (4k)
frame_vm_group_bin_21121 = frame (4k)
frame_vm_group_bin_21122 = frame (4k)
frame_vm_group_bin_21123 = frame (4k)
frame_vm_group_bin_21124 = frame (4k)
frame_vm_group_bin_21125 = frame (4k)
frame_vm_group_bin_21126 = frame (4k)
frame_vm_group_bin_21127 = frame (4k)
frame_vm_group_bin_21128 = frame (4k)
frame_vm_group_bin_21129 = frame (4k)
frame_vm_group_bin_2113 = frame (4k)
frame_vm_group_bin_21130 = frame (4k)
frame_vm_group_bin_21131 = frame (4k)
frame_vm_group_bin_21132 = frame (4k)
frame_vm_group_bin_21133 = frame (4k)
frame_vm_group_bin_21134 = frame (4k)
frame_vm_group_bin_21135 = frame (4k)
frame_vm_group_bin_21136 = frame (4k)
frame_vm_group_bin_21137 = frame (4k)
frame_vm_group_bin_21138 = frame (4k)
frame_vm_group_bin_21139 = frame (4k)
frame_vm_group_bin_2114 = frame (4k)
frame_vm_group_bin_21140 = frame (4k)
frame_vm_group_bin_21141 = frame (4k)
frame_vm_group_bin_21142 = frame (4k)
frame_vm_group_bin_21143 = frame (4k)
frame_vm_group_bin_21144 = frame (4k)
frame_vm_group_bin_21145 = frame (4k)
frame_vm_group_bin_21146 = frame (4k)
frame_vm_group_bin_21147 = frame (4k)
frame_vm_group_bin_21148 = frame (4k)
frame_vm_group_bin_21149 = frame (4k)
frame_vm_group_bin_2115 = frame (4k)
frame_vm_group_bin_21150 = frame (4k)
frame_vm_group_bin_21151 = frame (4k)
frame_vm_group_bin_21152 = frame (4k)
frame_vm_group_bin_21153 = frame (4k)
frame_vm_group_bin_21154 = frame (4k)
frame_vm_group_bin_21155 = frame (4k)
frame_vm_group_bin_21156 = frame (4k)
frame_vm_group_bin_21157 = frame (4k)
frame_vm_group_bin_21158 = frame (4k)
frame_vm_group_bin_21159 = frame (4k)
frame_vm_group_bin_2116 = frame (4k)
frame_vm_group_bin_21160 = frame (4k)
frame_vm_group_bin_21161 = frame (4k)
frame_vm_group_bin_21162 = frame (4k)
frame_vm_group_bin_21163 = frame (4k)
frame_vm_group_bin_21164 = frame (4k)
frame_vm_group_bin_21165 = frame (4k)
frame_vm_group_bin_21166 = frame (4k)
frame_vm_group_bin_21167 = frame (4k)
frame_vm_group_bin_21168 = frame (4k)
frame_vm_group_bin_21169 = frame (4k)
frame_vm_group_bin_2117 = frame (4k)
frame_vm_group_bin_21170 = frame (4k)
frame_vm_group_bin_21171 = frame (4k)
frame_vm_group_bin_21172 = frame (4k)
frame_vm_group_bin_21173 = frame (4k)
frame_vm_group_bin_21174 = frame (4k)
frame_vm_group_bin_21175 = frame (4k)
frame_vm_group_bin_21176 = frame (4k)
frame_vm_group_bin_21177 = frame (4k)
frame_vm_group_bin_21178 = frame (4k)
frame_vm_group_bin_21179 = frame (4k)
frame_vm_group_bin_2118 = frame (4k)
frame_vm_group_bin_21180 = frame (4k)
frame_vm_group_bin_21181 = frame (4k)
frame_vm_group_bin_21182 = frame (4k)
frame_vm_group_bin_21183 = frame (4k)
frame_vm_group_bin_21184 = frame (4k)
frame_vm_group_bin_21185 = frame (4k)
frame_vm_group_bin_21186 = frame (4k)
frame_vm_group_bin_21187 = frame (4k)
frame_vm_group_bin_21188 = frame (4k)
frame_vm_group_bin_21189 = frame (4k)
frame_vm_group_bin_2119 = frame (4k)
frame_vm_group_bin_21190 = frame (4k)
frame_vm_group_bin_21191 = frame (4k)
frame_vm_group_bin_21192 = frame (4k)
frame_vm_group_bin_21193 = frame (4k)
frame_vm_group_bin_21194 = frame (4k)
frame_vm_group_bin_21195 = frame (4k)
frame_vm_group_bin_21196 = frame (4k)
frame_vm_group_bin_21197 = frame (4k)
frame_vm_group_bin_21198 = frame (4k)
frame_vm_group_bin_21199 = frame (4k)
frame_vm_group_bin_2120 = frame (4k)
frame_vm_group_bin_21200 = frame (4k)
frame_vm_group_bin_21201 = frame (4k)
frame_vm_group_bin_21202 = frame (4k)
frame_vm_group_bin_21203 = frame (4k)
frame_vm_group_bin_21204 = frame (4k)
frame_vm_group_bin_21205 = frame (4k)
frame_vm_group_bin_21206 = frame (4k)
frame_vm_group_bin_21207 = frame (4k)
frame_vm_group_bin_21208 = frame (4k)
frame_vm_group_bin_21209 = frame (4k)
frame_vm_group_bin_2121 = frame (4k)
frame_vm_group_bin_21210 = frame (4k)
frame_vm_group_bin_21211 = frame (4k)
frame_vm_group_bin_21212 = frame (4k)
frame_vm_group_bin_21213 = frame (4k)
frame_vm_group_bin_21214 = frame (4k)
frame_vm_group_bin_21215 = frame (4k)
frame_vm_group_bin_21216 = frame (4k)
frame_vm_group_bin_21217 = frame (4k)
frame_vm_group_bin_21218 = frame (4k)
frame_vm_group_bin_21219 = frame (4k)
frame_vm_group_bin_2122 = frame (4k)
frame_vm_group_bin_21220 = frame (4k)
frame_vm_group_bin_21221 = frame (4k)
frame_vm_group_bin_21222 = frame (4k)
frame_vm_group_bin_21223 = frame (4k)
frame_vm_group_bin_21224 = frame (4k)
frame_vm_group_bin_21225 = frame (4k)
frame_vm_group_bin_21226 = frame (4k)
frame_vm_group_bin_21227 = frame (4k)
frame_vm_group_bin_21228 = frame (4k)
frame_vm_group_bin_21229 = frame (4k)
frame_vm_group_bin_2123 = frame (4k)
frame_vm_group_bin_21230 = frame (4k)
frame_vm_group_bin_21231 = frame (4k)
frame_vm_group_bin_21232 = frame (4k)
frame_vm_group_bin_21233 = frame (4k)
frame_vm_group_bin_21234 = frame (4k)
frame_vm_group_bin_21235 = frame (4k)
frame_vm_group_bin_21236 = frame (4k)
frame_vm_group_bin_21237 = frame (4k)
frame_vm_group_bin_21238 = frame (4k)
frame_vm_group_bin_21239 = frame (4k)
frame_vm_group_bin_2124 = frame (4k)
frame_vm_group_bin_21240 = frame (4k)
frame_vm_group_bin_21241 = frame (4k)
frame_vm_group_bin_21242 = frame (4k)
frame_vm_group_bin_21243 = frame (4k)
frame_vm_group_bin_21244 = frame (4k)
frame_vm_group_bin_21245 = frame (4k)
frame_vm_group_bin_21246 = frame (4k)
frame_vm_group_bin_21247 = frame (4k)
frame_vm_group_bin_21248 = frame (4k)
frame_vm_group_bin_21249 = frame (4k)
frame_vm_group_bin_2125 = frame (4k)
frame_vm_group_bin_21250 = frame (4k)
frame_vm_group_bin_21251 = frame (4k)
frame_vm_group_bin_21252 = frame (4k)
frame_vm_group_bin_21253 = frame (4k)
frame_vm_group_bin_21254 = frame (4k)
frame_vm_group_bin_21255 = frame (4k)
frame_vm_group_bin_21256 = frame (4k)
frame_vm_group_bin_21257 = frame (4k)
frame_vm_group_bin_21258 = frame (4k)
frame_vm_group_bin_21259 = frame (4k)
frame_vm_group_bin_2126 = frame (4k)
frame_vm_group_bin_21260 = frame (4k)
frame_vm_group_bin_21261 = frame (4k)
frame_vm_group_bin_21262 = frame (4k)
frame_vm_group_bin_21263 = frame (4k)
frame_vm_group_bin_21264 = frame (4k)
frame_vm_group_bin_21265 = frame (4k)
frame_vm_group_bin_21266 = frame (4k)
frame_vm_group_bin_21267 = frame (4k)
frame_vm_group_bin_21268 = frame (4k)
frame_vm_group_bin_21269 = frame (4k)
frame_vm_group_bin_2127 = frame (4k)
frame_vm_group_bin_21270 = frame (4k)
frame_vm_group_bin_21271 = frame (4k)
frame_vm_group_bin_21272 = frame (4k)
frame_vm_group_bin_21273 = frame (4k)
frame_vm_group_bin_21274 = frame (4k)
frame_vm_group_bin_21275 = frame (4k)
frame_vm_group_bin_21276 = frame (4k)
frame_vm_group_bin_21277 = frame (4k)
frame_vm_group_bin_21278 = frame (4k)
frame_vm_group_bin_21279 = frame (4k)
frame_vm_group_bin_2128 = frame (4k)
frame_vm_group_bin_21280 = frame (4k)
frame_vm_group_bin_21281 = frame (4k)
frame_vm_group_bin_21282 = frame (4k)
frame_vm_group_bin_21283 = frame (4k)
frame_vm_group_bin_21284 = frame (4k)
frame_vm_group_bin_21285 = frame (4k)
frame_vm_group_bin_21286 = frame (4k)
frame_vm_group_bin_21287 = frame (4k)
frame_vm_group_bin_21288 = frame (4k)
frame_vm_group_bin_21289 = frame (4k)
frame_vm_group_bin_2129 = frame (4k)
frame_vm_group_bin_21290 = frame (4k)
frame_vm_group_bin_21291 = frame (4k)
frame_vm_group_bin_21292 = frame (4k)
frame_vm_group_bin_21293 = frame (4k)
frame_vm_group_bin_21294 = frame (4k)
frame_vm_group_bin_21295 = frame (4k)
frame_vm_group_bin_21296 = frame (4k)
frame_vm_group_bin_21297 = frame (4k)
frame_vm_group_bin_21298 = frame (4k)
frame_vm_group_bin_21299 = frame (4k)
frame_vm_group_bin_2130 = frame (4k)
frame_vm_group_bin_21300 = frame (4k)
frame_vm_group_bin_21301 = frame (4k)
frame_vm_group_bin_21302 = frame (4k)
frame_vm_group_bin_21303 = frame (4k)
frame_vm_group_bin_21304 = frame (4k)
frame_vm_group_bin_21305 = frame (4k)
frame_vm_group_bin_21306 = frame (4k)
frame_vm_group_bin_21307 = frame (4k)
frame_vm_group_bin_21308 = frame (4k)
frame_vm_group_bin_21309 = frame (4k)
frame_vm_group_bin_2131 = frame (4k)
frame_vm_group_bin_21310 = frame (4k)
frame_vm_group_bin_21311 = frame (4k)
frame_vm_group_bin_21312 = frame (4k)
frame_vm_group_bin_21313 = frame (4k)
frame_vm_group_bin_21314 = frame (4k)
frame_vm_group_bin_21315 = frame (4k)
frame_vm_group_bin_21316 = frame (4k)
frame_vm_group_bin_21317 = frame (4k)
frame_vm_group_bin_21318 = frame (4k)
frame_vm_group_bin_21319 = frame (4k)
frame_vm_group_bin_2132 = frame (4k)
frame_vm_group_bin_21320 = frame (4k)
frame_vm_group_bin_21321 = frame (4k)
frame_vm_group_bin_21322 = frame (4k)
frame_vm_group_bin_21323 = frame (4k)
frame_vm_group_bin_21324 = frame (4k)
frame_vm_group_bin_21325 = frame (4k)
frame_vm_group_bin_21326 = frame (4k)
frame_vm_group_bin_21327 = frame (4k)
frame_vm_group_bin_21328 = frame (4k)
frame_vm_group_bin_21329 = frame (4k)
frame_vm_group_bin_2133 = frame (4k)
frame_vm_group_bin_21330 = frame (4k)
frame_vm_group_bin_21331 = frame (4k)
frame_vm_group_bin_21332 = frame (4k)
frame_vm_group_bin_21333 = frame (4k)
frame_vm_group_bin_21334 = frame (4k)
frame_vm_group_bin_21335 = frame (4k)
frame_vm_group_bin_21336 = frame (4k)
frame_vm_group_bin_21337 = frame (4k)
frame_vm_group_bin_21338 = frame (4k)
frame_vm_group_bin_21339 = frame (4k)
frame_vm_group_bin_2134 = frame (4k)
frame_vm_group_bin_21340 = frame (4k)
frame_vm_group_bin_21341 = frame (4k)
frame_vm_group_bin_21342 = frame (4k)
frame_vm_group_bin_21343 = frame (4k)
frame_vm_group_bin_21344 = frame (4k)
frame_vm_group_bin_21345 = frame (4k)
frame_vm_group_bin_21346 = frame (4k)
frame_vm_group_bin_21347 = frame (4k)
frame_vm_group_bin_21348 = frame (4k)
frame_vm_group_bin_21349 = frame (4k)
frame_vm_group_bin_2135 = frame (4k)
frame_vm_group_bin_21350 = frame (4k)
frame_vm_group_bin_21351 = frame (4k)
frame_vm_group_bin_21352 = frame (4k)
frame_vm_group_bin_21353 = frame (4k)
frame_vm_group_bin_21354 = frame (4k)
frame_vm_group_bin_21355 = frame (4k)
frame_vm_group_bin_21356 = frame (4k)
frame_vm_group_bin_21358 = frame (4k)
frame_vm_group_bin_21359 = frame (4k)
frame_vm_group_bin_2136 = frame (4k)
frame_vm_group_bin_21360 = frame (4k)
frame_vm_group_bin_21361 = frame (4k)
frame_vm_group_bin_21362 = frame (4k)
frame_vm_group_bin_21363 = frame (4k)
frame_vm_group_bin_21364 = frame (4k)
frame_vm_group_bin_21365 = frame (4k)
frame_vm_group_bin_21366 = frame (4k)
frame_vm_group_bin_21367 = frame (4k)
frame_vm_group_bin_21368 = frame (4k)
frame_vm_group_bin_21369 = frame (4k)
frame_vm_group_bin_2137 = frame (4k)
frame_vm_group_bin_21370 = frame (4k)
frame_vm_group_bin_21371 = frame (4k)
frame_vm_group_bin_21372 = frame (4k)
frame_vm_group_bin_21373 = frame (4k)
frame_vm_group_bin_21374 = frame (4k)
frame_vm_group_bin_21375 = frame (4k)
frame_vm_group_bin_21376 = frame (4k)
frame_vm_group_bin_21377 = frame (4k)
frame_vm_group_bin_21378 = frame (4k)
frame_vm_group_bin_21379 = frame (4k)
frame_vm_group_bin_2138 = frame (4k)
frame_vm_group_bin_21380 = frame (4k)
frame_vm_group_bin_21381 = frame (4k)
frame_vm_group_bin_21382 = frame (4k)
frame_vm_group_bin_21383 = frame (4k)
frame_vm_group_bin_21384 = frame (4k)
frame_vm_group_bin_21385 = frame (4k)
frame_vm_group_bin_21386 = frame (4k)
frame_vm_group_bin_21387 = frame (4k)
frame_vm_group_bin_21388 = frame (4k)
frame_vm_group_bin_21389 = frame (4k)
frame_vm_group_bin_2139 = frame (4k)
frame_vm_group_bin_21391 = frame (4k)
frame_vm_group_bin_21392 = frame (4k)
frame_vm_group_bin_21393 = frame (4k)
frame_vm_group_bin_21394 = frame (4k)
frame_vm_group_bin_21395 = frame (4k)
frame_vm_group_bin_21396 = frame (4k)
frame_vm_group_bin_21397 = frame (4k)
frame_vm_group_bin_21398 = frame (4k)
frame_vm_group_bin_21399 = frame (4k)
frame_vm_group_bin_2140 = frame (4k)
frame_vm_group_bin_21400 = frame (4k)
frame_vm_group_bin_21401 = frame (4k)
frame_vm_group_bin_21402 = frame (4k)
frame_vm_group_bin_21403 = frame (4k)
frame_vm_group_bin_21404 = frame (4k)
frame_vm_group_bin_21405 = frame (4k)
frame_vm_group_bin_21406 = frame (4k)
frame_vm_group_bin_21407 = frame (4k)
frame_vm_group_bin_21408 = frame (4k)
frame_vm_group_bin_21409 = frame (4k)
frame_vm_group_bin_2141 = frame (4k)
frame_vm_group_bin_21410 = frame (4k)
frame_vm_group_bin_21411 = frame (4k)
frame_vm_group_bin_21412 = frame (4k)
frame_vm_group_bin_21413 = frame (4k)
frame_vm_group_bin_21414 = frame (4k)
frame_vm_group_bin_21415 = frame (4k)
frame_vm_group_bin_21416 = frame (4k)
frame_vm_group_bin_21417 = frame (4k)
frame_vm_group_bin_21418 = frame (4k)
frame_vm_group_bin_21419 = frame (4k)
frame_vm_group_bin_2142 = frame (4k)
frame_vm_group_bin_21420 = frame (4k)
frame_vm_group_bin_21421 = frame (4k)
frame_vm_group_bin_21422 = frame (4k)
frame_vm_group_bin_21423 = frame (4k)
frame_vm_group_bin_21424 = frame (4k)
frame_vm_group_bin_21425 = frame (4k)
frame_vm_group_bin_21426 = frame (4k)
frame_vm_group_bin_21427 = frame (4k)
frame_vm_group_bin_21428 = frame (4k)
frame_vm_group_bin_21429 = frame (4k)
frame_vm_group_bin_2143 = frame (4k)
frame_vm_group_bin_21430 = frame (4k)
frame_vm_group_bin_21431 = frame (4k)
frame_vm_group_bin_21432 = frame (4k)
frame_vm_group_bin_21433 = frame (4k)
frame_vm_group_bin_21434 = frame (4k)
frame_vm_group_bin_21435 = frame (4k)
frame_vm_group_bin_21436 = frame (4k)
frame_vm_group_bin_21437 = frame (4k)
frame_vm_group_bin_21438 = frame (4k)
frame_vm_group_bin_21439 = frame (4k)
frame_vm_group_bin_2144 = frame (4k)
frame_vm_group_bin_21440 = frame (4k)
frame_vm_group_bin_21441 = frame (4k)
frame_vm_group_bin_21442 = frame (4k)
frame_vm_group_bin_21443 = frame (4k)
frame_vm_group_bin_21444 = frame (4k)
frame_vm_group_bin_21445 = frame (4k)
frame_vm_group_bin_21446 = frame (4k)
frame_vm_group_bin_21447 = frame (4k)
frame_vm_group_bin_21448 = frame (4k)
frame_vm_group_bin_21449 = frame (4k)
frame_vm_group_bin_2145 = frame (4k)
frame_vm_group_bin_21450 = frame (4k)
frame_vm_group_bin_21451 = frame (4k)
frame_vm_group_bin_21452 = frame (4k)
frame_vm_group_bin_21453 = frame (4k)
frame_vm_group_bin_21454 = frame (4k)
frame_vm_group_bin_21455 = frame (4k)
frame_vm_group_bin_21456 = frame (4k)
frame_vm_group_bin_21457 = frame (4k)
frame_vm_group_bin_21458 = frame (4k)
frame_vm_group_bin_21459 = frame (4k)
frame_vm_group_bin_2146 = frame (4k)
frame_vm_group_bin_21460 = frame (4k)
frame_vm_group_bin_21461 = frame (4k)
frame_vm_group_bin_21462 = frame (4k)
frame_vm_group_bin_21463 = frame (4k)
frame_vm_group_bin_21464 = frame (4k)
frame_vm_group_bin_21465 = frame (4k)
frame_vm_group_bin_21466 = frame (4k)
frame_vm_group_bin_21467 = frame (4k)
frame_vm_group_bin_21468 = frame (4k)
frame_vm_group_bin_21469 = frame (4k)
frame_vm_group_bin_2147 = frame (4k)
frame_vm_group_bin_21470 = frame (4k)
frame_vm_group_bin_21471 = frame (4k)
frame_vm_group_bin_21472 = frame (4k)
frame_vm_group_bin_21473 = frame (4k)
frame_vm_group_bin_21474 = frame (4k)
frame_vm_group_bin_21475 = frame (4k)
frame_vm_group_bin_21476 = frame (4k)
frame_vm_group_bin_21477 = frame (4k)
frame_vm_group_bin_21478 = frame (4k)
frame_vm_group_bin_21479 = frame (4k)
frame_vm_group_bin_2148 = frame (4k)
frame_vm_group_bin_21480 = frame (4k)
frame_vm_group_bin_21481 = frame (4k)
frame_vm_group_bin_21482 = frame (4k)
frame_vm_group_bin_21483 = frame (4k)
frame_vm_group_bin_21484 = frame (4k)
frame_vm_group_bin_21485 = frame (4k)
frame_vm_group_bin_21486 = frame (4k)
frame_vm_group_bin_21487 = frame (4k)
frame_vm_group_bin_21488 = frame (4k)
frame_vm_group_bin_21489 = frame (4k)
frame_vm_group_bin_2149 = frame (4k)
frame_vm_group_bin_21490 = frame (4k)
frame_vm_group_bin_21491 = frame (4k)
frame_vm_group_bin_21492 = frame (4k)
frame_vm_group_bin_21493 = frame (4k)
frame_vm_group_bin_21494 = frame (4k)
frame_vm_group_bin_21495 = frame (4k)
frame_vm_group_bin_21496 = frame (4k)
frame_vm_group_bin_21497 = frame (4k)
frame_vm_group_bin_21498 = frame (4k)
frame_vm_group_bin_21499 = frame (4k)
frame_vm_group_bin_2150 = frame (4k)
frame_vm_group_bin_21500 = frame (4k)
frame_vm_group_bin_21501 = frame (4k)
frame_vm_group_bin_21502 = frame (4k)
frame_vm_group_bin_21503 = frame (4k)
frame_vm_group_bin_21504 = frame (4k)
frame_vm_group_bin_21505 = frame (4k)
frame_vm_group_bin_21506 = frame (4k)
frame_vm_group_bin_21507 = frame (4k)
frame_vm_group_bin_21508 = frame (4k)
frame_vm_group_bin_21509 = frame (4k)
frame_vm_group_bin_2151 = frame (4k)
frame_vm_group_bin_21510 = frame (4k)
frame_vm_group_bin_21511 = frame (4k)
frame_vm_group_bin_21512 = frame (4k)
frame_vm_group_bin_21513 = frame (4k)
frame_vm_group_bin_21514 = frame (4k)
frame_vm_group_bin_21515 = frame (4k)
frame_vm_group_bin_21516 = frame (4k)
frame_vm_group_bin_21517 = frame (4k)
frame_vm_group_bin_21518 = frame (4k)
frame_vm_group_bin_21519 = frame (4k)
frame_vm_group_bin_2152 = frame (4k)
frame_vm_group_bin_21520 = frame (4k)
frame_vm_group_bin_21521 = frame (4k)
frame_vm_group_bin_21522 = frame (4k)
frame_vm_group_bin_21523 = frame (4k)
frame_vm_group_bin_21524 = frame (4k)
frame_vm_group_bin_21525 = frame (4k)
frame_vm_group_bin_21526 = frame (4k)
frame_vm_group_bin_21527 = frame (4k)
frame_vm_group_bin_21528 = frame (4k)
frame_vm_group_bin_21529 = frame (4k)
frame_vm_group_bin_2153 = frame (4k)
frame_vm_group_bin_21530 = frame (4k)
frame_vm_group_bin_21531 = frame (4k)
frame_vm_group_bin_21532 = frame (4k)
frame_vm_group_bin_21533 = frame (4k)
frame_vm_group_bin_21534 = frame (4k)
frame_vm_group_bin_21535 = frame (4k)
frame_vm_group_bin_21536 = frame (4k)
frame_vm_group_bin_21537 = frame (4k)
frame_vm_group_bin_21538 = frame (4k)
frame_vm_group_bin_21539 = frame (4k)
frame_vm_group_bin_2154 = frame (4k)
frame_vm_group_bin_21540 = frame (4k)
frame_vm_group_bin_21541 = frame (4k)
frame_vm_group_bin_21542 = frame (4k)
frame_vm_group_bin_21543 = frame (4k)
frame_vm_group_bin_21544 = frame (4k)
frame_vm_group_bin_21545 = frame (4k)
frame_vm_group_bin_21546 = frame (4k)
frame_vm_group_bin_21547 = frame (4k)
frame_vm_group_bin_21548 = frame (4k)
frame_vm_group_bin_21549 = frame (4k)
frame_vm_group_bin_2155 = frame (4k)
frame_vm_group_bin_21550 = frame (4k)
frame_vm_group_bin_21551 = frame (4k)
frame_vm_group_bin_21552 = frame (4k)
frame_vm_group_bin_21553 = frame (4k)
frame_vm_group_bin_21554 = frame (4k)
frame_vm_group_bin_21555 = frame (4k)
frame_vm_group_bin_21556 = frame (4k)
frame_vm_group_bin_21557 = frame (4k)
frame_vm_group_bin_21558 = frame (4k)
frame_vm_group_bin_21559 = frame (4k)
frame_vm_group_bin_2156 = frame (4k)
frame_vm_group_bin_21560 = frame (4k)
frame_vm_group_bin_21561 = frame (4k)
frame_vm_group_bin_21562 = frame (4k)
frame_vm_group_bin_21563 = frame (4k)
frame_vm_group_bin_21564 = frame (4k)
frame_vm_group_bin_21565 = frame (4k)
frame_vm_group_bin_21566 = frame (4k)
frame_vm_group_bin_21567 = frame (4k)
frame_vm_group_bin_21568 = frame (4k)
frame_vm_group_bin_21569 = frame (4k)
frame_vm_group_bin_2157 = frame (4k)
frame_vm_group_bin_21570 = frame (4k)
frame_vm_group_bin_21571 = frame (4k)
frame_vm_group_bin_21572 = frame (4k)
frame_vm_group_bin_21573 = frame (4k)
frame_vm_group_bin_21574 = frame (4k)
frame_vm_group_bin_21575 = frame (4k)
frame_vm_group_bin_21576 = frame (4k)
frame_vm_group_bin_21577 = frame (4k)
frame_vm_group_bin_21578 = frame (4k)
frame_vm_group_bin_21579 = frame (4k)
frame_vm_group_bin_2158 = frame (4k)
frame_vm_group_bin_21580 = frame (4k)
frame_vm_group_bin_21581 = frame (4k)
frame_vm_group_bin_21582 = frame (4k)
frame_vm_group_bin_21583 = frame (4k)
frame_vm_group_bin_21584 = frame (4k)
frame_vm_group_bin_21585 = frame (4k)
frame_vm_group_bin_21586 = frame (4k)
frame_vm_group_bin_21587 = frame (4k)
frame_vm_group_bin_21588 = frame (4k)
frame_vm_group_bin_21589 = frame (4k)
frame_vm_group_bin_2159 = frame (4k)
frame_vm_group_bin_21590 = frame (4k)
frame_vm_group_bin_21591 = frame (4k)
frame_vm_group_bin_21592 = frame (4k)
frame_vm_group_bin_21593 = frame (4k)
frame_vm_group_bin_21594 = frame (4k)
frame_vm_group_bin_21595 = frame (4k)
frame_vm_group_bin_21596 = frame (4k)
frame_vm_group_bin_21597 = frame (4k)
frame_vm_group_bin_21598 = frame (4k)
frame_vm_group_bin_21599 = frame (4k)
frame_vm_group_bin_2160 = frame (4k)
frame_vm_group_bin_21600 = frame (4k)
frame_vm_group_bin_21601 = frame (4k)
frame_vm_group_bin_21602 = frame (4k)
frame_vm_group_bin_21603 = frame (4k)
frame_vm_group_bin_21604 = frame (4k)
frame_vm_group_bin_21605 = frame (4k)
frame_vm_group_bin_21606 = frame (4k)
frame_vm_group_bin_21607 = frame (4k)
frame_vm_group_bin_21608 = frame (4k)
frame_vm_group_bin_21609 = frame (4k)
frame_vm_group_bin_2161 = frame (4k)
frame_vm_group_bin_21610 = frame (4k)
frame_vm_group_bin_21611 = frame (4k)
frame_vm_group_bin_21612 = frame (4k)
frame_vm_group_bin_21613 = frame (4k)
frame_vm_group_bin_21614 = frame (4k)
frame_vm_group_bin_21615 = frame (4k)
frame_vm_group_bin_21616 = frame (4k)
frame_vm_group_bin_21617 = frame (4k)
frame_vm_group_bin_21618 = frame (4k)
frame_vm_group_bin_21619 = frame (4k)
frame_vm_group_bin_2162 = frame (4k)
frame_vm_group_bin_21620 = frame (4k)
frame_vm_group_bin_21621 = frame (4k)
frame_vm_group_bin_21622 = frame (4k)
frame_vm_group_bin_21623 = frame (4k)
frame_vm_group_bin_21624 = frame (4k)
frame_vm_group_bin_21625 = frame (4k)
frame_vm_group_bin_21626 = frame (4k)
frame_vm_group_bin_21627 = frame (4k)
frame_vm_group_bin_21628 = frame (4k)
frame_vm_group_bin_21629 = frame (4k)
frame_vm_group_bin_2163 = frame (4k)
frame_vm_group_bin_21630 = frame (4k)
frame_vm_group_bin_21631 = frame (4k)
frame_vm_group_bin_21632 = frame (4k)
frame_vm_group_bin_21633 = frame (4k)
frame_vm_group_bin_21634 = frame (4k)
frame_vm_group_bin_21635 = frame (4k)
frame_vm_group_bin_21636 = frame (4k)
frame_vm_group_bin_21637 = frame (4k)
frame_vm_group_bin_21638 = frame (4k)
frame_vm_group_bin_21639 = frame (4k)
frame_vm_group_bin_2164 = frame (4k)
frame_vm_group_bin_21640 = frame (4k)
frame_vm_group_bin_21641 = frame (4k)
frame_vm_group_bin_21642 = frame (4k)
frame_vm_group_bin_21643 = frame (4k)
frame_vm_group_bin_21644 = frame (4k)
frame_vm_group_bin_21645 = frame (4k)
frame_vm_group_bin_21646 = frame (4k)
frame_vm_group_bin_21647 = frame (4k)
frame_vm_group_bin_21648 = frame (4k)
frame_vm_group_bin_21649 = frame (4k)
frame_vm_group_bin_2165 = frame (4k)
frame_vm_group_bin_21650 = frame (4k)
frame_vm_group_bin_21651 = frame (4k)
frame_vm_group_bin_21652 = frame (4k)
frame_vm_group_bin_21653 = frame (4k)
frame_vm_group_bin_21654 = frame (4k)
frame_vm_group_bin_21655 = frame (4k)
frame_vm_group_bin_21656 = frame (4k)
frame_vm_group_bin_21657 = frame (4k)
frame_vm_group_bin_21658 = frame (4k)
frame_vm_group_bin_21659 = frame (4k)
frame_vm_group_bin_2166 = frame (4k)
frame_vm_group_bin_21660 = frame (4k)
frame_vm_group_bin_21661 = frame (4k)
frame_vm_group_bin_21662 = frame (4k)
frame_vm_group_bin_21663 = frame (4k)
frame_vm_group_bin_21664 = frame (4k)
frame_vm_group_bin_21665 = frame (4k)
frame_vm_group_bin_21666 = frame (4k)
frame_vm_group_bin_21667 = frame (4k)
frame_vm_group_bin_21668 = frame (4k)
frame_vm_group_bin_21669 = frame (4k)
frame_vm_group_bin_2167 = frame (4k)
frame_vm_group_bin_21670 = frame (4k)
frame_vm_group_bin_21671 = frame (4k)
frame_vm_group_bin_21672 = frame (4k)
frame_vm_group_bin_21673 = frame (4k)
frame_vm_group_bin_21674 = frame (4k)
frame_vm_group_bin_21675 = frame (4k)
frame_vm_group_bin_21676 = frame (4k)
frame_vm_group_bin_21677 = frame (4k)
frame_vm_group_bin_21678 = frame (4k)
frame_vm_group_bin_21679 = frame (4k)
frame_vm_group_bin_2168 = frame (4k)
frame_vm_group_bin_21680 = frame (4k)
frame_vm_group_bin_21681 = frame (4k)
frame_vm_group_bin_21682 = frame (4k)
frame_vm_group_bin_21683 = frame (4k)
frame_vm_group_bin_21684 = frame (4k)
frame_vm_group_bin_21685 = frame (4k)
frame_vm_group_bin_21686 = frame (4k)
frame_vm_group_bin_21687 = frame (4k)
frame_vm_group_bin_21688 = frame (4k)
frame_vm_group_bin_21689 = frame (4k)
frame_vm_group_bin_2169 = frame (4k)
frame_vm_group_bin_21690 = frame (4k)
frame_vm_group_bin_21691 = frame (4k)
frame_vm_group_bin_21692 = frame (4k)
frame_vm_group_bin_21693 = frame (4k)
frame_vm_group_bin_21694 = frame (4k)
frame_vm_group_bin_21695 = frame (4k)
frame_vm_group_bin_21696 = frame (4k)
frame_vm_group_bin_21697 = frame (4k)
frame_vm_group_bin_21698 = frame (4k)
frame_vm_group_bin_21699 = frame (4k)
frame_vm_group_bin_2170 = frame (4k)
frame_vm_group_bin_21700 = frame (4k)
frame_vm_group_bin_21701 = frame (4k)
frame_vm_group_bin_21702 = frame (4k)
frame_vm_group_bin_21703 = frame (4k)
frame_vm_group_bin_21704 = frame (4k)
frame_vm_group_bin_21705 = frame (4k)
frame_vm_group_bin_21706 = frame (4k)
frame_vm_group_bin_21707 = frame (4k)
frame_vm_group_bin_21708 = frame (4k)
frame_vm_group_bin_21709 = frame (4k)
frame_vm_group_bin_2171 = frame (4k)
frame_vm_group_bin_21710 = frame (4k)
frame_vm_group_bin_21711 = frame (4k)
frame_vm_group_bin_21712 = frame (4k)
frame_vm_group_bin_21713 = frame (4k)
frame_vm_group_bin_21714 = frame (4k)
frame_vm_group_bin_21715 = frame (4k)
frame_vm_group_bin_21716 = frame (4k)
frame_vm_group_bin_21717 = frame (4k)
frame_vm_group_bin_21718 = frame (4k)
frame_vm_group_bin_21719 = frame (4k)
frame_vm_group_bin_2172 = frame (4k)
frame_vm_group_bin_21720 = frame (4k)
frame_vm_group_bin_21721 = frame (4k)
frame_vm_group_bin_21722 = frame (4k)
frame_vm_group_bin_21723 = frame (4k)
frame_vm_group_bin_21724 = frame (4k)
frame_vm_group_bin_21725 = frame (4k)
frame_vm_group_bin_21726 = frame (4k)
frame_vm_group_bin_21727 = frame (4k)
frame_vm_group_bin_21728 = frame (4k)
frame_vm_group_bin_21729 = frame (4k)
frame_vm_group_bin_2173 = frame (4k)
frame_vm_group_bin_21730 = frame (4k)
frame_vm_group_bin_21731 = frame (4k)
frame_vm_group_bin_21732 = frame (4k)
frame_vm_group_bin_21733 = frame (4k)
frame_vm_group_bin_21734 = frame (4k)
frame_vm_group_bin_21735 = frame (4k)
frame_vm_group_bin_21736 = frame (4k)
frame_vm_group_bin_21737 = frame (4k)
frame_vm_group_bin_21738 = frame (4k)
frame_vm_group_bin_21739 = frame (4k)
frame_vm_group_bin_2174 = frame (4k)
frame_vm_group_bin_21740 = frame (4k)
frame_vm_group_bin_21741 = frame (4k)
frame_vm_group_bin_21742 = frame (4k)
frame_vm_group_bin_21743 = frame (4k)
frame_vm_group_bin_21744 = frame (4k)
frame_vm_group_bin_21745 = frame (4k)
frame_vm_group_bin_21746 = frame (4k)
frame_vm_group_bin_21747 = frame (4k)
frame_vm_group_bin_21748 = frame (4k)
frame_vm_group_bin_21749 = frame (4k)
frame_vm_group_bin_2175 = frame (4k)
frame_vm_group_bin_21750 = frame (4k)
frame_vm_group_bin_21751 = frame (4k)
frame_vm_group_bin_21752 = frame (4k)
frame_vm_group_bin_21753 = frame (4k)
frame_vm_group_bin_21754 = frame (4k)
frame_vm_group_bin_21755 = frame (4k)
frame_vm_group_bin_21756 = frame (4k)
frame_vm_group_bin_21757 = frame (4k)
frame_vm_group_bin_21758 = frame (4k)
frame_vm_group_bin_21759 = frame (4k)
frame_vm_group_bin_2176 = frame (4k)
frame_vm_group_bin_21760 = frame (4k)
frame_vm_group_bin_21761 = frame (4k)
frame_vm_group_bin_21762 = frame (4k)
frame_vm_group_bin_21763 = frame (4k)
frame_vm_group_bin_21764 = frame (4k)
frame_vm_group_bin_21765 = frame (4k)
frame_vm_group_bin_21766 = frame (4k)
frame_vm_group_bin_21767 = frame (4k)
frame_vm_group_bin_21768 = frame (4k)
frame_vm_group_bin_21769 = frame (4k)
frame_vm_group_bin_2177 = frame (4k)
frame_vm_group_bin_21770 = frame (4k)
frame_vm_group_bin_21771 = frame (4k)
frame_vm_group_bin_21772 = frame (4k)
frame_vm_group_bin_21773 = frame (4k)
frame_vm_group_bin_21774 = frame (4k)
frame_vm_group_bin_21775 = frame (4k)
frame_vm_group_bin_21776 = frame (4k)
frame_vm_group_bin_21777 = frame (4k)
frame_vm_group_bin_21778 = frame (4k)
frame_vm_group_bin_21779 = frame (4k)
frame_vm_group_bin_2178 = frame (4k)
frame_vm_group_bin_21780 = frame (4k)
frame_vm_group_bin_21781 = frame (4k)
frame_vm_group_bin_21782 = frame (4k)
frame_vm_group_bin_21783 = frame (4k)
frame_vm_group_bin_21784 = frame (4k)
frame_vm_group_bin_21785 = frame (4k)
frame_vm_group_bin_21786 = frame (4k)
frame_vm_group_bin_21787 = frame (4k)
frame_vm_group_bin_21788 = frame (4k)
frame_vm_group_bin_21789 = frame (4k)
frame_vm_group_bin_2179 = frame (4k)
frame_vm_group_bin_21790 = frame (4k)
frame_vm_group_bin_21791 = frame (4k)
frame_vm_group_bin_21792 = frame (4k)
frame_vm_group_bin_21793 = frame (4k)
frame_vm_group_bin_21794 = frame (4k)
frame_vm_group_bin_21795 = frame (4k)
frame_vm_group_bin_21796 = frame (4k)
frame_vm_group_bin_21797 = frame (4k)
frame_vm_group_bin_21798 = frame (4k)
frame_vm_group_bin_21799 = frame (4k)
frame_vm_group_bin_2180 = frame (4k)
frame_vm_group_bin_21800 = frame (4k)
frame_vm_group_bin_21801 = frame (4k)
frame_vm_group_bin_21802 = frame (4k)
frame_vm_group_bin_21803 = frame (4k)
frame_vm_group_bin_21804 = frame (4k)
frame_vm_group_bin_21805 = frame (4k)
frame_vm_group_bin_21806 = frame (4k)
frame_vm_group_bin_21807 = frame (4k)
frame_vm_group_bin_21808 = frame (4k)
frame_vm_group_bin_21809 = frame (4k)
frame_vm_group_bin_2181 = frame (4k)
frame_vm_group_bin_21810 = frame (4k)
frame_vm_group_bin_21811 = frame (4k)
frame_vm_group_bin_21812 = frame (4k)
frame_vm_group_bin_21813 = frame (4k)
frame_vm_group_bin_21814 = frame (4k)
frame_vm_group_bin_21815 = frame (4k)
frame_vm_group_bin_21816 = frame (4k)
frame_vm_group_bin_21817 = frame (4k)
frame_vm_group_bin_21818 = frame (4k)
frame_vm_group_bin_21819 = frame (4k)
frame_vm_group_bin_2182 = frame (4k)
frame_vm_group_bin_21820 = frame (4k)
frame_vm_group_bin_21821 = frame (4k)
frame_vm_group_bin_21822 = frame (4k)
frame_vm_group_bin_21823 = frame (4k)
frame_vm_group_bin_21824 = frame (4k)
frame_vm_group_bin_21825 = frame (4k)
frame_vm_group_bin_21826 = frame (4k)
frame_vm_group_bin_21827 = frame (4k)
frame_vm_group_bin_21828 = frame (4k)
frame_vm_group_bin_21829 = frame (4k)
frame_vm_group_bin_2183 = frame (4k)
frame_vm_group_bin_21830 = frame (4k)
frame_vm_group_bin_21831 = frame (4k)
frame_vm_group_bin_21832 = frame (4k)
frame_vm_group_bin_21833 = frame (4k)
frame_vm_group_bin_21834 = frame (4k)
frame_vm_group_bin_21835 = frame (4k)
frame_vm_group_bin_21836 = frame (4k)
frame_vm_group_bin_21837 = frame (4k)
frame_vm_group_bin_21838 = frame (4k)
frame_vm_group_bin_21839 = frame (4k)
frame_vm_group_bin_2184 = frame (4k)
frame_vm_group_bin_21840 = frame (4k)
frame_vm_group_bin_21841 = frame (4k)
frame_vm_group_bin_21842 = frame (4k)
frame_vm_group_bin_21843 = frame (4k)
frame_vm_group_bin_21844 = frame (4k)
frame_vm_group_bin_21845 = frame (4k)
frame_vm_group_bin_21846 = frame (4k)
frame_vm_group_bin_21847 = frame (4k)
frame_vm_group_bin_21848 = frame (4k)
frame_vm_group_bin_21849 = frame (4k)
frame_vm_group_bin_2185 = frame (4k)
frame_vm_group_bin_21850 = frame (4k)
frame_vm_group_bin_21851 = frame (4k)
frame_vm_group_bin_21852 = frame (4k)
frame_vm_group_bin_21853 = frame (4k)
frame_vm_group_bin_21854 = frame (4k)
frame_vm_group_bin_21855 = frame (4k)
frame_vm_group_bin_21856 = frame (4k)
frame_vm_group_bin_21857 = frame (4k)
frame_vm_group_bin_21858 = frame (4k)
frame_vm_group_bin_21859 = frame (4k)
frame_vm_group_bin_2186 = frame (4k)
frame_vm_group_bin_21860 = frame (4k)
frame_vm_group_bin_21861 = frame (4k)
frame_vm_group_bin_21862 = frame (4k)
frame_vm_group_bin_21863 = frame (4k)
frame_vm_group_bin_21864 = frame (4k)
frame_vm_group_bin_21865 = frame (4k)
frame_vm_group_bin_21866 = frame (4k)
frame_vm_group_bin_21867 = frame (4k)
frame_vm_group_bin_21868 = frame (4k)
frame_vm_group_bin_21869 = frame (4k)
frame_vm_group_bin_2187 = frame (4k)
frame_vm_group_bin_21870 = frame (4k)
frame_vm_group_bin_21871 = frame (4k)
frame_vm_group_bin_21872 = frame (4k)
frame_vm_group_bin_21873 = frame (4k)
frame_vm_group_bin_21874 = frame (4k)
frame_vm_group_bin_21875 = frame (4k)
frame_vm_group_bin_21876 = frame (4k)
frame_vm_group_bin_21877 = frame (4k)
frame_vm_group_bin_21878 = frame (4k)
frame_vm_group_bin_21879 = frame (4k)
frame_vm_group_bin_2188 = frame (4k)
frame_vm_group_bin_21880 = frame (4k)
frame_vm_group_bin_21881 = frame (4k)
frame_vm_group_bin_21882 = frame (4k)
frame_vm_group_bin_21883 = frame (4k)
frame_vm_group_bin_21884 = frame (4k)
frame_vm_group_bin_21885 = frame (4k)
frame_vm_group_bin_21886 = frame (4k)
frame_vm_group_bin_21887 = frame (4k)
frame_vm_group_bin_21888 = frame (4k)
frame_vm_group_bin_21889 = frame (4k)
frame_vm_group_bin_2189 = frame (4k)
frame_vm_group_bin_21890 = frame (4k)
frame_vm_group_bin_21891 = frame (4k)
frame_vm_group_bin_21892 = frame (4k)
frame_vm_group_bin_21893 = frame (4k)
frame_vm_group_bin_21894 = frame (4k)
frame_vm_group_bin_21895 = frame (4k)
frame_vm_group_bin_21896 = frame (4k)
frame_vm_group_bin_21897 = frame (4k)
frame_vm_group_bin_21898 = frame (4k)
frame_vm_group_bin_21899 = frame (4k)
frame_vm_group_bin_2190 = frame (4k)
frame_vm_group_bin_21900 = frame (4k)
frame_vm_group_bin_21901 = frame (4k)
frame_vm_group_bin_21902 = frame (4k)
frame_vm_group_bin_21903 = frame (4k)
frame_vm_group_bin_21904 = frame (4k)
frame_vm_group_bin_21905 = frame (4k)
frame_vm_group_bin_21906 = frame (4k)
frame_vm_group_bin_21907 = frame (4k)
frame_vm_group_bin_21908 = frame (4k)
frame_vm_group_bin_21909 = frame (4k)
frame_vm_group_bin_2191 = frame (4k)
frame_vm_group_bin_21910 = frame (4k)
frame_vm_group_bin_21911 = frame (4k)
frame_vm_group_bin_21912 = frame (4k)
frame_vm_group_bin_21913 = frame (4k)
frame_vm_group_bin_21914 = frame (4k)
frame_vm_group_bin_21915 = frame (4k)
frame_vm_group_bin_21916 = frame (4k)
frame_vm_group_bin_21917 = frame (4k)
frame_vm_group_bin_21918 = frame (4k)
frame_vm_group_bin_21919 = frame (4k)
frame_vm_group_bin_2192 = frame (4k)
frame_vm_group_bin_21920 = frame (4k)
frame_vm_group_bin_21921 = frame (4k)
frame_vm_group_bin_21922 = frame (4k)
frame_vm_group_bin_21923 = frame (4k)
frame_vm_group_bin_21924 = frame (4k)
frame_vm_group_bin_21925 = frame (4k)
frame_vm_group_bin_21926 = frame (4k)
frame_vm_group_bin_21927 = frame (4k)
frame_vm_group_bin_21928 = frame (4k)
frame_vm_group_bin_21929 = frame (4k)
frame_vm_group_bin_2193 = frame (4k)
frame_vm_group_bin_21930 = frame (4k)
frame_vm_group_bin_21931 = frame (4k)
frame_vm_group_bin_21932 = frame (4k)
frame_vm_group_bin_21933 = frame (4k)
frame_vm_group_bin_21934 = frame (4k)
frame_vm_group_bin_21935 = frame (4k)
frame_vm_group_bin_21936 = frame (4k)
frame_vm_group_bin_21937 = frame (4k)
frame_vm_group_bin_21938 = frame (4k)
frame_vm_group_bin_21939 = frame (4k)
frame_vm_group_bin_2194 = frame (4k)
frame_vm_group_bin_21940 = frame (4k)
frame_vm_group_bin_21941 = frame (4k)
frame_vm_group_bin_21942 = frame (4k)
frame_vm_group_bin_21943 = frame (4k)
frame_vm_group_bin_21944 = frame (4k)
frame_vm_group_bin_21945 = frame (4k)
frame_vm_group_bin_21946 = frame (4k)
frame_vm_group_bin_21947 = frame (4k)
frame_vm_group_bin_21948 = frame (4k)
frame_vm_group_bin_21949 = frame (4k)
frame_vm_group_bin_2195 = frame (4k)
frame_vm_group_bin_21950 = frame (4k)
frame_vm_group_bin_21951 = frame (4k)
frame_vm_group_bin_21952 = frame (4k)
frame_vm_group_bin_21953 = frame (4k)
frame_vm_group_bin_21954 = frame (4k)
frame_vm_group_bin_21955 = frame (4k)
frame_vm_group_bin_21956 = frame (4k)
frame_vm_group_bin_21957 = frame (4k)
frame_vm_group_bin_21958 = frame (4k)
frame_vm_group_bin_21959 = frame (4k)
frame_vm_group_bin_2196 = frame (4k)
frame_vm_group_bin_21960 = frame (4k)
frame_vm_group_bin_21961 = frame (4k)
frame_vm_group_bin_21962 = frame (4k)
frame_vm_group_bin_21963 = frame (4k)
frame_vm_group_bin_21964 = frame (4k)
frame_vm_group_bin_21965 = frame (4k)
frame_vm_group_bin_21966 = frame (4k)
frame_vm_group_bin_21967 = frame (4k)
frame_vm_group_bin_21968 = frame (4k)
frame_vm_group_bin_21969 = frame (4k)
frame_vm_group_bin_2197 = frame (4k)
frame_vm_group_bin_21970 = frame (4k)
frame_vm_group_bin_21971 = frame (4k)
frame_vm_group_bin_21972 = frame (4k)
frame_vm_group_bin_21973 = frame (4k)
frame_vm_group_bin_21974 = frame (4k)
frame_vm_group_bin_21975 = frame (4k)
frame_vm_group_bin_21976 = frame (4k)
frame_vm_group_bin_21977 = frame (4k)
frame_vm_group_bin_21978 = frame (4k)
frame_vm_group_bin_21979 = frame (4k)
frame_vm_group_bin_2198 = frame (4k)
frame_vm_group_bin_21980 = frame (4k)
frame_vm_group_bin_21981 = frame (4k)
frame_vm_group_bin_21982 = frame (4k)
frame_vm_group_bin_21983 = frame (4k)
frame_vm_group_bin_21984 = frame (4k)
frame_vm_group_bin_21985 = frame (4k)
frame_vm_group_bin_21986 = frame (4k)
frame_vm_group_bin_21987 = frame (4k)
frame_vm_group_bin_21988 = frame (4k)
frame_vm_group_bin_21989 = frame (4k)
frame_vm_group_bin_2199 = frame (4k)
frame_vm_group_bin_21990 = frame (4k)
frame_vm_group_bin_21991 = frame (4k)
frame_vm_group_bin_21992 = frame (4k)
frame_vm_group_bin_21993 = frame (4k)
frame_vm_group_bin_21994 = frame (4k)
frame_vm_group_bin_21995 = frame (4k)
frame_vm_group_bin_21996 = frame (4k)
frame_vm_group_bin_21997 = frame (4k)
frame_vm_group_bin_21998 = frame (4k)
frame_vm_group_bin_21999 = frame (4k)
frame_vm_group_bin_2200 = frame (4k)
frame_vm_group_bin_22000 = frame (4k)
frame_vm_group_bin_22001 = frame (4k)
frame_vm_group_bin_22002 = frame (4k)
frame_vm_group_bin_22003 = frame (4k)
frame_vm_group_bin_22004 = frame (4k)
frame_vm_group_bin_22005 = frame (4k)
frame_vm_group_bin_22006 = frame (4k)
frame_vm_group_bin_22007 = frame (4k)
frame_vm_group_bin_22008 = frame (4k)
frame_vm_group_bin_22009 = frame (4k)
frame_vm_group_bin_2201 = frame (4k)
frame_vm_group_bin_22010 = frame (4k)
frame_vm_group_bin_22011 = frame (4k)
frame_vm_group_bin_22012 = frame (4k)
frame_vm_group_bin_22013 = frame (4k)
frame_vm_group_bin_22014 = frame (4k)
frame_vm_group_bin_22015 = frame (4k)
frame_vm_group_bin_22016 = frame (4k)
frame_vm_group_bin_22017 = frame (4k)
frame_vm_group_bin_22018 = frame (4k)
frame_vm_group_bin_22019 = frame (4k)
frame_vm_group_bin_2202 = frame (4k)
frame_vm_group_bin_22020 = frame (4k)
frame_vm_group_bin_22021 = frame (4k)
frame_vm_group_bin_22022 = frame (4k)
frame_vm_group_bin_22023 = frame (4k)
frame_vm_group_bin_22024 = frame (4k)
frame_vm_group_bin_22025 = frame (4k)
frame_vm_group_bin_22026 = frame (4k)
frame_vm_group_bin_22027 = frame (4k)
frame_vm_group_bin_22028 = frame (4k)
frame_vm_group_bin_22029 = frame (4k)
frame_vm_group_bin_2203 = frame (4k)
frame_vm_group_bin_22030 = frame (4k)
frame_vm_group_bin_22031 = frame (4k)
frame_vm_group_bin_22032 = frame (4k)
frame_vm_group_bin_22033 = frame (4k)
frame_vm_group_bin_22034 = frame (4k)
frame_vm_group_bin_22035 = frame (4k)
frame_vm_group_bin_22036 = frame (4k)
frame_vm_group_bin_22037 = frame (4k)
frame_vm_group_bin_22038 = frame (4k)
frame_vm_group_bin_22039 = frame (4k)
frame_vm_group_bin_2204 = frame (4k)
frame_vm_group_bin_22040 = frame (4k)
frame_vm_group_bin_22041 = frame (4k)
frame_vm_group_bin_22042 = frame (4k)
frame_vm_group_bin_22043 = frame (4k)
frame_vm_group_bin_22044 = frame (4k)
frame_vm_group_bin_22045 = frame (4k)
frame_vm_group_bin_22046 = frame (4k)
frame_vm_group_bin_22047 = frame (4k)
frame_vm_group_bin_22048 = frame (4k)
frame_vm_group_bin_22049 = frame (4k)
frame_vm_group_bin_2205 = frame (4k)
frame_vm_group_bin_22050 = frame (4k)
frame_vm_group_bin_22051 = frame (4k)
frame_vm_group_bin_22052 = frame (4k)
frame_vm_group_bin_22053 = frame (4k)
frame_vm_group_bin_22054 = frame (4k)
frame_vm_group_bin_22055 = frame (4k)
frame_vm_group_bin_22056 = frame (4k)
frame_vm_group_bin_22057 = frame (4k)
frame_vm_group_bin_22058 = frame (4k)
frame_vm_group_bin_22059 = frame (4k)
frame_vm_group_bin_2206 = frame (4k)
frame_vm_group_bin_22060 = frame (4k)
frame_vm_group_bin_22061 = frame (4k)
frame_vm_group_bin_22062 = frame (4k)
frame_vm_group_bin_22063 = frame (4k)
frame_vm_group_bin_22064 = frame (4k)
frame_vm_group_bin_22065 = frame (4k)
frame_vm_group_bin_22066 = frame (4k)
frame_vm_group_bin_22067 = frame (4k)
frame_vm_group_bin_22068 = frame (4k)
frame_vm_group_bin_22069 = frame (4k)
frame_vm_group_bin_2207 = frame (4k)
frame_vm_group_bin_22070 = frame (4k)
frame_vm_group_bin_22071 = frame (4k)
frame_vm_group_bin_22072 = frame (4k)
frame_vm_group_bin_22073 = frame (4k)
frame_vm_group_bin_22074 = frame (4k)
frame_vm_group_bin_22075 = frame (4k)
frame_vm_group_bin_22076 = frame (4k)
frame_vm_group_bin_22077 = frame (4k)
frame_vm_group_bin_22078 = frame (4k)
frame_vm_group_bin_22079 = frame (4k)
frame_vm_group_bin_2208 = frame (4k)
frame_vm_group_bin_22080 = frame (4k)
frame_vm_group_bin_22081 = frame (4k)
frame_vm_group_bin_22082 = frame (4k)
frame_vm_group_bin_22083 = frame (4k)
frame_vm_group_bin_22084 = frame (4k)
frame_vm_group_bin_22085 = frame (4k)
frame_vm_group_bin_22086 = frame (4k)
frame_vm_group_bin_22087 = frame (4k)
frame_vm_group_bin_22088 = frame (4k)
frame_vm_group_bin_22089 = frame (4k)
frame_vm_group_bin_2209 = frame (4k)
frame_vm_group_bin_22090 = frame (4k)
frame_vm_group_bin_22091 = frame (4k)
frame_vm_group_bin_22092 = frame (4k)
frame_vm_group_bin_22093 = frame (4k)
frame_vm_group_bin_22094 = frame (4k)
frame_vm_group_bin_22095 = frame (4k)
frame_vm_group_bin_22096 = frame (4k)
frame_vm_group_bin_22097 = frame (4k)
frame_vm_group_bin_22098 = frame (4k)
frame_vm_group_bin_22099 = frame (4k)
frame_vm_group_bin_2210 = frame (4k)
frame_vm_group_bin_22100 = frame (4k)
frame_vm_group_bin_22101 = frame (4k)
frame_vm_group_bin_22102 = frame (4k)
frame_vm_group_bin_22103 = frame (4k)
frame_vm_group_bin_22104 = frame (4k)
frame_vm_group_bin_22105 = frame (4k)
frame_vm_group_bin_22106 = frame (4k)
frame_vm_group_bin_22107 = frame (4k)
frame_vm_group_bin_22108 = frame (4k)
frame_vm_group_bin_22109 = frame (4k)
frame_vm_group_bin_2211 = frame (4k)
frame_vm_group_bin_22110 = frame (4k)
frame_vm_group_bin_22111 = frame (4k)
frame_vm_group_bin_22112 = frame (4k)
frame_vm_group_bin_22113 = frame (4k)
frame_vm_group_bin_22114 = frame (4k)
frame_vm_group_bin_22115 = frame (4k)
frame_vm_group_bin_22116 = frame (4k)
frame_vm_group_bin_22117 = frame (4k)
frame_vm_group_bin_22118 = frame (4k)
frame_vm_group_bin_22119 = frame (4k)
frame_vm_group_bin_2212 = frame (4k)
frame_vm_group_bin_22120 = frame (4k)
frame_vm_group_bin_22121 = frame (4k)
frame_vm_group_bin_22122 = frame (4k)
frame_vm_group_bin_22123 = frame (4k)
frame_vm_group_bin_22124 = frame (4k)
frame_vm_group_bin_22125 = frame (4k)
frame_vm_group_bin_22126 = frame (4k)
frame_vm_group_bin_22127 = frame (4k)
frame_vm_group_bin_22128 = frame (4k)
frame_vm_group_bin_22129 = frame (4k)
frame_vm_group_bin_2213 = frame (4k)
frame_vm_group_bin_22130 = frame (4k)
frame_vm_group_bin_22131 = frame (4k)
frame_vm_group_bin_22132 = frame (4k)
frame_vm_group_bin_22133 = frame (4k)
frame_vm_group_bin_22134 = frame (4k)
frame_vm_group_bin_22135 = frame (4k)
frame_vm_group_bin_22136 = frame (4k)
frame_vm_group_bin_22137 = frame (4k)
frame_vm_group_bin_22138 = frame (4k)
frame_vm_group_bin_22139 = frame (4k)
frame_vm_group_bin_2214 = frame (4k)
frame_vm_group_bin_22140 = frame (4k)
frame_vm_group_bin_22141 = frame (4k)
frame_vm_group_bin_22142 = frame (4k)
frame_vm_group_bin_22143 = frame (4k)
frame_vm_group_bin_22144 = frame (4k)
frame_vm_group_bin_22145 = frame (4k)
frame_vm_group_bin_22146 = frame (4k)
frame_vm_group_bin_22147 = frame (4k)
frame_vm_group_bin_22148 = frame (4k)
frame_vm_group_bin_22149 = frame (4k)
frame_vm_group_bin_2215 = frame (4k)
frame_vm_group_bin_22150 = frame (4k)
frame_vm_group_bin_22151 = frame (4k)
frame_vm_group_bin_22152 = frame (4k)
frame_vm_group_bin_22153 = frame (4k)
frame_vm_group_bin_22154 = frame (4k)
frame_vm_group_bin_22155 = frame (4k)
frame_vm_group_bin_22156 = frame (4k)
frame_vm_group_bin_22157 = frame (4k)
frame_vm_group_bin_22158 = frame (4k)
frame_vm_group_bin_22159 = frame (4k)
frame_vm_group_bin_2216 = frame (4k)
frame_vm_group_bin_22160 = frame (4k)
frame_vm_group_bin_22161 = frame (4k)
frame_vm_group_bin_22162 = frame (4k)
frame_vm_group_bin_22163 = frame (4k)
frame_vm_group_bin_22164 = frame (4k)
frame_vm_group_bin_22165 = frame (4k)
frame_vm_group_bin_22166 = frame (4k)
frame_vm_group_bin_22167 = frame (4k)
frame_vm_group_bin_22168 = frame (4k)
frame_vm_group_bin_22169 = frame (4k)
frame_vm_group_bin_2217 = frame (4k)
frame_vm_group_bin_22170 = frame (4k)
frame_vm_group_bin_22171 = frame (4k)
frame_vm_group_bin_22172 = frame (4k)
frame_vm_group_bin_22173 = frame (4k)
frame_vm_group_bin_22174 = frame (4k)
frame_vm_group_bin_22175 = frame (4k)
frame_vm_group_bin_22176 = frame (4k)
frame_vm_group_bin_22177 = frame (4k)
frame_vm_group_bin_22178 = frame (4k)
frame_vm_group_bin_22179 = frame (4k)
frame_vm_group_bin_2218 = frame (4k)
frame_vm_group_bin_22180 = frame (4k)
frame_vm_group_bin_22181 = frame (4k)
frame_vm_group_bin_22182 = frame (4k)
frame_vm_group_bin_22183 = frame (4k)
frame_vm_group_bin_22184 = frame (4k)
frame_vm_group_bin_22185 = frame (4k)
frame_vm_group_bin_22186 = frame (4k)
frame_vm_group_bin_22187 = frame (4k)
frame_vm_group_bin_22188 = frame (4k)
frame_vm_group_bin_22189 = frame (4k)
frame_vm_group_bin_2219 = frame (4k)
frame_vm_group_bin_22190 = frame (4k)
frame_vm_group_bin_22191 = frame (4k)
frame_vm_group_bin_22192 = frame (4k)
frame_vm_group_bin_22193 = frame (4k)
frame_vm_group_bin_22194 = frame (4k)
frame_vm_group_bin_22195 = frame (4k)
frame_vm_group_bin_22196 = frame (4k)
frame_vm_group_bin_22197 = frame (4k)
frame_vm_group_bin_22198 = frame (4k)
frame_vm_group_bin_22199 = frame (4k)
frame_vm_group_bin_2220 = frame (4k)
frame_vm_group_bin_22200 = frame (4k)
frame_vm_group_bin_22201 = frame (4k)
frame_vm_group_bin_22202 = frame (4k)
frame_vm_group_bin_22203 = frame (4k)
frame_vm_group_bin_22204 = frame (4k)
frame_vm_group_bin_22205 = frame (4k)
frame_vm_group_bin_22206 = frame (4k)
frame_vm_group_bin_22207 = frame (4k)
frame_vm_group_bin_22208 = frame (4k)
frame_vm_group_bin_22209 = frame (4k)
frame_vm_group_bin_2221 = frame (4k)
frame_vm_group_bin_22210 = frame (4k)
frame_vm_group_bin_22211 = frame (4k)
frame_vm_group_bin_22212 = frame (4k)
frame_vm_group_bin_22213 = frame (4k)
frame_vm_group_bin_22214 = frame (4k)
frame_vm_group_bin_22215 = frame (4k)
frame_vm_group_bin_22216 = frame (4k)
frame_vm_group_bin_22217 = frame (4k)
frame_vm_group_bin_22218 = frame (4k)
frame_vm_group_bin_22219 = frame (4k)
frame_vm_group_bin_2222 = frame (4k)
frame_vm_group_bin_22220 = frame (4k)
frame_vm_group_bin_22221 = frame (4k)
frame_vm_group_bin_22222 = frame (4k)
frame_vm_group_bin_22223 = frame (4k)
frame_vm_group_bin_22224 = frame (4k)
frame_vm_group_bin_22225 = frame (4k)
frame_vm_group_bin_22226 = frame (4k)
frame_vm_group_bin_22227 = frame (4k)
frame_vm_group_bin_22228 = frame (4k)
frame_vm_group_bin_22229 = frame (4k)
frame_vm_group_bin_2223 = frame (4k)
frame_vm_group_bin_22230 = frame (4k)
frame_vm_group_bin_22231 = frame (4k)
frame_vm_group_bin_22232 = frame (4k)
frame_vm_group_bin_22233 = frame (4k)
frame_vm_group_bin_22234 = frame (4k)
frame_vm_group_bin_22235 = frame (4k)
frame_vm_group_bin_22236 = frame (4k)
frame_vm_group_bin_22237 = frame (4k)
frame_vm_group_bin_22238 = frame (4k)
frame_vm_group_bin_22239 = frame (4k)
frame_vm_group_bin_2224 = frame (4k)
frame_vm_group_bin_22240 = frame (4k)
frame_vm_group_bin_22241 = frame (4k)
frame_vm_group_bin_22242 = frame (4k)
frame_vm_group_bin_22243 = frame (4k)
frame_vm_group_bin_22244 = frame (4k)
frame_vm_group_bin_22245 = frame (4k)
frame_vm_group_bin_22246 = frame (4k)
frame_vm_group_bin_22247 = frame (4k)
frame_vm_group_bin_22248 = frame (4k)
frame_vm_group_bin_22249 = frame (4k)
frame_vm_group_bin_2225 = frame (4k)
frame_vm_group_bin_22250 = frame (4k)
frame_vm_group_bin_22251 = frame (4k)
frame_vm_group_bin_22252 = frame (4k)
frame_vm_group_bin_22253 = frame (4k)
frame_vm_group_bin_22254 = frame (4k)
frame_vm_group_bin_22255 = frame (4k)
frame_vm_group_bin_22256 = frame (4k)
frame_vm_group_bin_22257 = frame (4k)
frame_vm_group_bin_22258 = frame (4k)
frame_vm_group_bin_22259 = frame (4k)
frame_vm_group_bin_2226 = frame (4k)
frame_vm_group_bin_22260 = frame (4k)
frame_vm_group_bin_22261 = frame (4k)
frame_vm_group_bin_22262 = frame (4k)
frame_vm_group_bin_22263 = frame (4k)
frame_vm_group_bin_22264 = frame (4k)
frame_vm_group_bin_22265 = frame (4k)
frame_vm_group_bin_22266 = frame (4k)
frame_vm_group_bin_22267 = frame (4k)
frame_vm_group_bin_22268 = frame (4k)
frame_vm_group_bin_22269 = frame (4k)
frame_vm_group_bin_2227 = frame (4k)
frame_vm_group_bin_22270 = frame (4k)
frame_vm_group_bin_22271 = frame (4k)
frame_vm_group_bin_22272 = frame (4k)
frame_vm_group_bin_22273 = frame (4k)
frame_vm_group_bin_22274 = frame (4k)
frame_vm_group_bin_22275 = frame (4k)
frame_vm_group_bin_22276 = frame (4k)
frame_vm_group_bin_22277 = frame (4k)
frame_vm_group_bin_22278 = frame (4k)
frame_vm_group_bin_22279 = frame (4k)
frame_vm_group_bin_2228 = frame (4k)
frame_vm_group_bin_22280 = frame (4k)
frame_vm_group_bin_22281 = frame (4k)
frame_vm_group_bin_22282 = frame (4k)
frame_vm_group_bin_22283 = frame (4k)
frame_vm_group_bin_22284 = frame (4k)
frame_vm_group_bin_22285 = frame (4k)
frame_vm_group_bin_22286 = frame (4k)
frame_vm_group_bin_22287 = frame (4k)
frame_vm_group_bin_22288 = frame (4k)
frame_vm_group_bin_22289 = frame (4k)
frame_vm_group_bin_2229 = frame (4k)
frame_vm_group_bin_22290 = frame (4k)
frame_vm_group_bin_22291 = frame (4k)
frame_vm_group_bin_22292 = frame (4k)
frame_vm_group_bin_22293 = frame (4k)
frame_vm_group_bin_22294 = frame (4k)
frame_vm_group_bin_22295 = frame (4k)
frame_vm_group_bin_22296 = frame (4k)
frame_vm_group_bin_22297 = frame (4k)
frame_vm_group_bin_22298 = frame (4k)
frame_vm_group_bin_22299 = frame (4k)
frame_vm_group_bin_2230 = frame (4k)
frame_vm_group_bin_22300 = frame (4k)
frame_vm_group_bin_22301 = frame (4k)
frame_vm_group_bin_22302 = frame (4k)
frame_vm_group_bin_22303 = frame (4k)
frame_vm_group_bin_22304 = frame (4k)
frame_vm_group_bin_22305 = frame (4k)
frame_vm_group_bin_22306 = frame (4k)
frame_vm_group_bin_22307 = frame (4k)
frame_vm_group_bin_22308 = frame (4k)
frame_vm_group_bin_22309 = frame (4k)
frame_vm_group_bin_2231 = frame (4k)
frame_vm_group_bin_22310 = frame (4k)
frame_vm_group_bin_22311 = frame (4k)
frame_vm_group_bin_22312 = frame (4k)
frame_vm_group_bin_22313 = frame (4k)
frame_vm_group_bin_22314 = frame (4k)
frame_vm_group_bin_22315 = frame (4k)
frame_vm_group_bin_22316 = frame (4k)
frame_vm_group_bin_22317 = frame (4k)
frame_vm_group_bin_22318 = frame (4k)
frame_vm_group_bin_22319 = frame (4k)
frame_vm_group_bin_2232 = frame (4k)
frame_vm_group_bin_22320 = frame (4k)
frame_vm_group_bin_22321 = frame (4k)
frame_vm_group_bin_22322 = frame (4k)
frame_vm_group_bin_22323 = frame (4k)
frame_vm_group_bin_22324 = frame (4k)
frame_vm_group_bin_22325 = frame (4k)
frame_vm_group_bin_22326 = frame (4k)
frame_vm_group_bin_22327 = frame (4k)
frame_vm_group_bin_22328 = frame (4k)
frame_vm_group_bin_22329 = frame (4k)
frame_vm_group_bin_2233 = frame (4k)
frame_vm_group_bin_22330 = frame (4k)
frame_vm_group_bin_22331 = frame (4k)
frame_vm_group_bin_22332 = frame (4k)
frame_vm_group_bin_22333 = frame (4k)
frame_vm_group_bin_22334 = frame (4k)
frame_vm_group_bin_22335 = frame (4k)
frame_vm_group_bin_22336 = frame (4k)
frame_vm_group_bin_22337 = frame (4k)
frame_vm_group_bin_22338 = frame (4k)
frame_vm_group_bin_22339 = frame (4k)
frame_vm_group_bin_2234 = frame (4k)
frame_vm_group_bin_22340 = frame (4k)
frame_vm_group_bin_22341 = frame (4k)
frame_vm_group_bin_22342 = frame (4k)
frame_vm_group_bin_22343 = frame (4k)
frame_vm_group_bin_22344 = frame (4k)
frame_vm_group_bin_22345 = frame (4k)
frame_vm_group_bin_22346 = frame (4k)
frame_vm_group_bin_22347 = frame (4k)
frame_vm_group_bin_22348 = frame (4k)
frame_vm_group_bin_22349 = frame (4k)
frame_vm_group_bin_2235 = frame (4k)
frame_vm_group_bin_22350 = frame (4k)
frame_vm_group_bin_22351 = frame (4k)
frame_vm_group_bin_22352 = frame (4k)
frame_vm_group_bin_22353 = frame (4k)
frame_vm_group_bin_22354 = frame (4k)
frame_vm_group_bin_22355 = frame (4k)
frame_vm_group_bin_22356 = frame (4k)
frame_vm_group_bin_22357 = frame (4k)
frame_vm_group_bin_22358 = frame (4k)
frame_vm_group_bin_22359 = frame (4k)
frame_vm_group_bin_2236 = frame (4k)
frame_vm_group_bin_22360 = frame (4k)
frame_vm_group_bin_22361 = frame (4k)
frame_vm_group_bin_22362 = frame (4k)
frame_vm_group_bin_22363 = frame (4k)
frame_vm_group_bin_22364 = frame (4k)
frame_vm_group_bin_22365 = frame (4k)
frame_vm_group_bin_22366 = frame (4k)
frame_vm_group_bin_22367 = frame (4k)
frame_vm_group_bin_22368 = frame (4k)
frame_vm_group_bin_22369 = frame (4k)
frame_vm_group_bin_2237 = frame (4k)
frame_vm_group_bin_22370 = frame (4k)
frame_vm_group_bin_22371 = frame (4k)
frame_vm_group_bin_22372 = frame (4k)
frame_vm_group_bin_22373 = frame (4k)
frame_vm_group_bin_22374 = frame (4k)
frame_vm_group_bin_22375 = frame (4k)
frame_vm_group_bin_22376 = frame (4k)
frame_vm_group_bin_22377 = frame (4k)
frame_vm_group_bin_22378 = frame (4k)
frame_vm_group_bin_22379 = frame (4k)
frame_vm_group_bin_2238 = frame (4k)
frame_vm_group_bin_22380 = frame (4k)
frame_vm_group_bin_22381 = frame (4k)
frame_vm_group_bin_22382 = frame (4k)
frame_vm_group_bin_22383 = frame (4k)
frame_vm_group_bin_22384 = frame (4k)
frame_vm_group_bin_22385 = frame (4k)
frame_vm_group_bin_22386 = frame (4k)
frame_vm_group_bin_22387 = frame (4k)
frame_vm_group_bin_22388 = frame (4k)
frame_vm_group_bin_22389 = frame (4k)
frame_vm_group_bin_2239 = frame (4k)
frame_vm_group_bin_22390 = frame (4k)
frame_vm_group_bin_22391 = frame (4k)
frame_vm_group_bin_22392 = frame (4k)
frame_vm_group_bin_22393 = frame (4k)
frame_vm_group_bin_22394 = frame (4k)
frame_vm_group_bin_22395 = frame (4k)
frame_vm_group_bin_22396 = frame (4k)
frame_vm_group_bin_22397 = frame (4k)
frame_vm_group_bin_22398 = frame (4k)
frame_vm_group_bin_22399 = frame (4k)
frame_vm_group_bin_2240 = frame (4k)
frame_vm_group_bin_22400 = frame (4k)
frame_vm_group_bin_22401 = frame (4k)
frame_vm_group_bin_22402 = frame (4k)
frame_vm_group_bin_22403 = frame (4k)
frame_vm_group_bin_22404 = frame (4k)
frame_vm_group_bin_22405 = frame (4k)
frame_vm_group_bin_22406 = frame (4k)
frame_vm_group_bin_22407 = frame (4k)
frame_vm_group_bin_22408 = frame (4k)
frame_vm_group_bin_22409 = frame (4k)
frame_vm_group_bin_2241 = frame (4k)
frame_vm_group_bin_22410 = frame (4k)
frame_vm_group_bin_22411 = frame (4k)
frame_vm_group_bin_22412 = frame (4k)
frame_vm_group_bin_22413 = frame (4k)
frame_vm_group_bin_22414 = frame (4k)
frame_vm_group_bin_22415 = frame (4k)
frame_vm_group_bin_22416 = frame (4k)
frame_vm_group_bin_22417 = frame (4k)
frame_vm_group_bin_22418 = frame (4k)
frame_vm_group_bin_22419 = frame (4k)
frame_vm_group_bin_2242 = frame (4k)
frame_vm_group_bin_22420 = frame (4k)
frame_vm_group_bin_22421 = frame (4k)
frame_vm_group_bin_22422 = frame (4k)
frame_vm_group_bin_22423 = frame (4k)
frame_vm_group_bin_22424 = frame (4k)
frame_vm_group_bin_22425 = frame (4k)
frame_vm_group_bin_22426 = frame (4k)
frame_vm_group_bin_22427 = frame (4k)
frame_vm_group_bin_22428 = frame (4k)
frame_vm_group_bin_22429 = frame (4k)
frame_vm_group_bin_2243 = frame (4k)
frame_vm_group_bin_22430 = frame (4k)
frame_vm_group_bin_22431 = frame (4k)
frame_vm_group_bin_22432 = frame (4k)
frame_vm_group_bin_22433 = frame (4k)
frame_vm_group_bin_22434 = frame (4k)
frame_vm_group_bin_22435 = frame (4k)
frame_vm_group_bin_22436 = frame (4k)
frame_vm_group_bin_22437 = frame (4k)
frame_vm_group_bin_22438 = frame (4k)
frame_vm_group_bin_22439 = frame (4k)
frame_vm_group_bin_2244 = frame (4k)
frame_vm_group_bin_22440 = frame (4k)
frame_vm_group_bin_22441 = frame (4k)
frame_vm_group_bin_22442 = frame (4k)
frame_vm_group_bin_22443 = frame (4k)
frame_vm_group_bin_22444 = frame (4k)
frame_vm_group_bin_22445 = frame (4k)
frame_vm_group_bin_22446 = frame (4k)
frame_vm_group_bin_22447 = frame (4k)
frame_vm_group_bin_22448 = frame (4k)
frame_vm_group_bin_22449 = frame (4k)
frame_vm_group_bin_2245 = frame (4k)
frame_vm_group_bin_22450 = frame (4k)
frame_vm_group_bin_22451 = frame (4k)
frame_vm_group_bin_22452 = frame (4k)
frame_vm_group_bin_22453 = frame (4k)
frame_vm_group_bin_22454 = frame (4k)
frame_vm_group_bin_22455 = frame (4k)
frame_vm_group_bin_22456 = frame (4k)
frame_vm_group_bin_22457 = frame (4k)
frame_vm_group_bin_22458 = frame (4k)
frame_vm_group_bin_22459 = frame (4k)
frame_vm_group_bin_2246 = frame (4k)
frame_vm_group_bin_22460 = frame (4k)
frame_vm_group_bin_22461 = frame (4k)
frame_vm_group_bin_22462 = frame (4k)
frame_vm_group_bin_22463 = frame (4k)
frame_vm_group_bin_22464 = frame (4k)
frame_vm_group_bin_22465 = frame (4k)
frame_vm_group_bin_22466 = frame (4k)
frame_vm_group_bin_22467 = frame (4k)
frame_vm_group_bin_22468 = frame (4k)
frame_vm_group_bin_22469 = frame (4k)
frame_vm_group_bin_2247 = frame (4k)
frame_vm_group_bin_22470 = frame (4k)
frame_vm_group_bin_22471 = frame (4k)
frame_vm_group_bin_22472 = frame (4k)
frame_vm_group_bin_22473 = frame (4k)
frame_vm_group_bin_22474 = frame (4k)
frame_vm_group_bin_22475 = frame (4k)
frame_vm_group_bin_22476 = frame (4k)
frame_vm_group_bin_22477 = frame (4k)
frame_vm_group_bin_22478 = frame (4k)
frame_vm_group_bin_22479 = frame (4k)
frame_vm_group_bin_2248 = frame (4k)
frame_vm_group_bin_22480 = frame (4k)
frame_vm_group_bin_22481 = frame (4k)
frame_vm_group_bin_22482 = frame (4k)
frame_vm_group_bin_22483 = frame (4k)
frame_vm_group_bin_22484 = frame (4k)
frame_vm_group_bin_22485 = frame (4k)
frame_vm_group_bin_22486 = frame (4k)
frame_vm_group_bin_22487 = frame (4k)
frame_vm_group_bin_22488 = frame (4k)
frame_vm_group_bin_22489 = frame (4k)
frame_vm_group_bin_2249 = frame (4k)
frame_vm_group_bin_22490 = frame (4k)
frame_vm_group_bin_22491 = frame (4k)
frame_vm_group_bin_22492 = frame (4k)
frame_vm_group_bin_22493 = frame (4k)
frame_vm_group_bin_22494 = frame (4k)
frame_vm_group_bin_22495 = frame (4k)
frame_vm_group_bin_22496 = frame (4k)
frame_vm_group_bin_22497 = frame (4k)
frame_vm_group_bin_22498 = frame (4k)
frame_vm_group_bin_22499 = frame (4k)
frame_vm_group_bin_2250 = frame (4k)
frame_vm_group_bin_22500 = frame (4k)
frame_vm_group_bin_22501 = frame (4k)
frame_vm_group_bin_22502 = frame (4k)
frame_vm_group_bin_22503 = frame (4k)
frame_vm_group_bin_22504 = frame (4k)
frame_vm_group_bin_22505 = frame (4k)
frame_vm_group_bin_22506 = frame (4k)
frame_vm_group_bin_22507 = frame (4k)
frame_vm_group_bin_22508 = frame (4k)
frame_vm_group_bin_22509 = frame (4k)
frame_vm_group_bin_2251 = frame (4k)
frame_vm_group_bin_22510 = frame (4k)
frame_vm_group_bin_22511 = frame (4k)
frame_vm_group_bin_22512 = frame (4k)
frame_vm_group_bin_22513 = frame (4k)
frame_vm_group_bin_22514 = frame (4k)
frame_vm_group_bin_22515 = frame (4k)
frame_vm_group_bin_22516 = frame (4k)
frame_vm_group_bin_22517 = frame (4k)
frame_vm_group_bin_22518 = frame (4k)
frame_vm_group_bin_22519 = frame (4k)
frame_vm_group_bin_2252 = frame (4k)
frame_vm_group_bin_22520 = frame (4k)
frame_vm_group_bin_22521 = frame (4k)
frame_vm_group_bin_22522 = frame (4k)
frame_vm_group_bin_22523 = frame (4k)
frame_vm_group_bin_22524 = frame (4k)
frame_vm_group_bin_22525 = frame (4k)
frame_vm_group_bin_22526 = frame (4k)
frame_vm_group_bin_22527 = frame (4k)
frame_vm_group_bin_22528 = frame (4k)
frame_vm_group_bin_22529 = frame (4k)
frame_vm_group_bin_2253 = frame (4k)
frame_vm_group_bin_22530 = frame (4k)
frame_vm_group_bin_22531 = frame (4k)
frame_vm_group_bin_22532 = frame (4k)
frame_vm_group_bin_22533 = frame (4k)
frame_vm_group_bin_22534 = frame (4k)
frame_vm_group_bin_22535 = frame (4k)
frame_vm_group_bin_22536 = frame (4k)
frame_vm_group_bin_22537 = frame (4k)
frame_vm_group_bin_22538 = frame (4k)
frame_vm_group_bin_22539 = frame (4k)
frame_vm_group_bin_2254 = frame (4k)
frame_vm_group_bin_22540 = frame (4k)
frame_vm_group_bin_22541 = frame (4k)
frame_vm_group_bin_22542 = frame (4k)
frame_vm_group_bin_22543 = frame (4k)
frame_vm_group_bin_22544 = frame (4k)
frame_vm_group_bin_22545 = frame (4k)
frame_vm_group_bin_22546 = frame (4k)
frame_vm_group_bin_22547 = frame (4k)
frame_vm_group_bin_22548 = frame (4k)
frame_vm_group_bin_22549 = frame (4k)
frame_vm_group_bin_2255 = frame (4k)
frame_vm_group_bin_22550 = frame (4k)
frame_vm_group_bin_22551 = frame (4k)
frame_vm_group_bin_22552 = frame (4k)
frame_vm_group_bin_22553 = frame (4k)
frame_vm_group_bin_22554 = frame (4k)
frame_vm_group_bin_22555 = frame (4k)
frame_vm_group_bin_22556 = frame (4k)
frame_vm_group_bin_22557 = frame (4k)
frame_vm_group_bin_22558 = frame (4k)
frame_vm_group_bin_22559 = frame (4k)
frame_vm_group_bin_2256 = frame (4k)
frame_vm_group_bin_22560 = frame (4k)
frame_vm_group_bin_22561 = frame (4k)
frame_vm_group_bin_22562 = frame (4k)
frame_vm_group_bin_22563 = frame (4k)
frame_vm_group_bin_22564 = frame (4k)
frame_vm_group_bin_22565 = frame (4k)
frame_vm_group_bin_22566 = frame (4k)
frame_vm_group_bin_22567 = frame (4k)
frame_vm_group_bin_22568 = frame (4k)
frame_vm_group_bin_22569 = frame (4k)
frame_vm_group_bin_2257 = frame (4k)
frame_vm_group_bin_22570 = frame (4k)
frame_vm_group_bin_22571 = frame (4k)
frame_vm_group_bin_22572 = frame (4k)
frame_vm_group_bin_22573 = frame (4k)
frame_vm_group_bin_22574 = frame (4k)
frame_vm_group_bin_22575 = frame (4k)
frame_vm_group_bin_22576 = frame (4k)
frame_vm_group_bin_22577 = frame (4k)
frame_vm_group_bin_22578 = frame (4k)
frame_vm_group_bin_22579 = frame (4k)
frame_vm_group_bin_2258 = frame (4k)
frame_vm_group_bin_22580 = frame (4k)
frame_vm_group_bin_22581 = frame (4k)
frame_vm_group_bin_22582 = frame (4k)
frame_vm_group_bin_22583 = frame (4k)
frame_vm_group_bin_22584 = frame (4k)
frame_vm_group_bin_22585 = frame (4k)
frame_vm_group_bin_22586 = frame (4k)
frame_vm_group_bin_22587 = frame (4k)
frame_vm_group_bin_22588 = frame (4k)
frame_vm_group_bin_22589 = frame (4k)
frame_vm_group_bin_2259 = frame (4k)
frame_vm_group_bin_22590 = frame (4k)
frame_vm_group_bin_22591 = frame (4k)
frame_vm_group_bin_22592 = frame (4k)
frame_vm_group_bin_22593 = frame (4k)
frame_vm_group_bin_22594 = frame (4k)
frame_vm_group_bin_22595 = frame (4k)
frame_vm_group_bin_22596 = frame (4k)
frame_vm_group_bin_22597 = frame (4k)
frame_vm_group_bin_22598 = frame (4k)
frame_vm_group_bin_22599 = frame (4k)
frame_vm_group_bin_2260 = frame (4k)
frame_vm_group_bin_22600 = frame (4k)
frame_vm_group_bin_22601 = frame (4k)
frame_vm_group_bin_22602 = frame (4k)
frame_vm_group_bin_22603 = frame (4k)
frame_vm_group_bin_22604 = frame (4k)
frame_vm_group_bin_22605 = frame (4k)
frame_vm_group_bin_22606 = frame (4k)
frame_vm_group_bin_22607 = frame (4k)
frame_vm_group_bin_22608 = frame (4k)
frame_vm_group_bin_22609 = frame (4k)
frame_vm_group_bin_2261 = frame (4k)
frame_vm_group_bin_22610 = frame (4k)
frame_vm_group_bin_22611 = frame (4k)
frame_vm_group_bin_22612 = frame (4k)
frame_vm_group_bin_22613 = frame (4k)
frame_vm_group_bin_22614 = frame (4k)
frame_vm_group_bin_22615 = frame (4k)
frame_vm_group_bin_22616 = frame (4k)
frame_vm_group_bin_22617 = frame (4k)
frame_vm_group_bin_22618 = frame (4k)
frame_vm_group_bin_22619 = frame (4k)
frame_vm_group_bin_2262 = frame (4k)
frame_vm_group_bin_22620 = frame (4k)
frame_vm_group_bin_22621 = frame (4k)
frame_vm_group_bin_22622 = frame (4k)
frame_vm_group_bin_22623 = frame (4k)
frame_vm_group_bin_22624 = frame (4k)
frame_vm_group_bin_22625 = frame (4k)
frame_vm_group_bin_22626 = frame (4k)
frame_vm_group_bin_22627 = frame (4k)
frame_vm_group_bin_22628 = frame (4k)
frame_vm_group_bin_22629 = frame (4k)
frame_vm_group_bin_2263 = frame (4k)
frame_vm_group_bin_22630 = frame (4k)
frame_vm_group_bin_22631 = frame (4k)
frame_vm_group_bin_22632 = frame (4k)
frame_vm_group_bin_22633 = frame (4k)
frame_vm_group_bin_22634 = frame (4k)
frame_vm_group_bin_22635 = frame (4k)
frame_vm_group_bin_22636 = frame (4k)
frame_vm_group_bin_22637 = frame (4k)
frame_vm_group_bin_22638 = frame (4k)
frame_vm_group_bin_22639 = frame (4k)
frame_vm_group_bin_2264 = frame (4k)
frame_vm_group_bin_22640 = frame (4k)
frame_vm_group_bin_22641 = frame (4k)
frame_vm_group_bin_22642 = frame (4k)
frame_vm_group_bin_22643 = frame (4k)
frame_vm_group_bin_22644 = frame (4k)
frame_vm_group_bin_22645 = frame (4k)
frame_vm_group_bin_22646 = frame (4k)
frame_vm_group_bin_22647 = frame (4k)
frame_vm_group_bin_22648 = frame (4k)
frame_vm_group_bin_22649 = frame (4k)
frame_vm_group_bin_2265 = frame (4k)
frame_vm_group_bin_22650 = frame (4k)
frame_vm_group_bin_22651 = frame (4k)
frame_vm_group_bin_22652 = frame (4k)
frame_vm_group_bin_22653 = frame (4k)
frame_vm_group_bin_22654 = frame (4k)
frame_vm_group_bin_22655 = frame (4k)
frame_vm_group_bin_22656 = frame (4k)
frame_vm_group_bin_22657 = frame (4k)
frame_vm_group_bin_22658 = frame (4k)
frame_vm_group_bin_22659 = frame (4k)
frame_vm_group_bin_2266 = frame (4k)
frame_vm_group_bin_22660 = frame (4k)
frame_vm_group_bin_22661 = frame (4k)
frame_vm_group_bin_22662 = frame (4k)
frame_vm_group_bin_22663 = frame (4k)
frame_vm_group_bin_22664 = frame (4k)
frame_vm_group_bin_22665 = frame (4k)
frame_vm_group_bin_22666 = frame (4k)
frame_vm_group_bin_22667 = frame (4k)
frame_vm_group_bin_22668 = frame (4k)
frame_vm_group_bin_22669 = frame (4k)
frame_vm_group_bin_2267 = frame (4k)
frame_vm_group_bin_22670 = frame (4k)
frame_vm_group_bin_22671 = frame (4k)
frame_vm_group_bin_22672 = frame (4k)
frame_vm_group_bin_22673 = frame (4k)
frame_vm_group_bin_22674 = frame (4k)
frame_vm_group_bin_22675 = frame (4k)
frame_vm_group_bin_22676 = frame (4k)
frame_vm_group_bin_22677 = frame (4k)
frame_vm_group_bin_22678 = frame (4k)
frame_vm_group_bin_22679 = frame (4k)
frame_vm_group_bin_2268 = frame (4k)
frame_vm_group_bin_22680 = frame (4k)
frame_vm_group_bin_22681 = frame (4k)
frame_vm_group_bin_22682 = frame (4k)
frame_vm_group_bin_22683 = frame (4k)
frame_vm_group_bin_22684 = frame (4k)
frame_vm_group_bin_22685 = frame (4k)
frame_vm_group_bin_22686 = frame (4k)
frame_vm_group_bin_22687 = frame (4k)
frame_vm_group_bin_22688 = frame (4k)
frame_vm_group_bin_22689 = frame (4k)
frame_vm_group_bin_2269 = frame (4k)
frame_vm_group_bin_22690 = frame (4k)
frame_vm_group_bin_22691 = frame (4k)
frame_vm_group_bin_22692 = frame (4k)
frame_vm_group_bin_22693 = frame (4k)
frame_vm_group_bin_22694 = frame (4k)
frame_vm_group_bin_22695 = frame (4k)
frame_vm_group_bin_22696 = frame (4k)
frame_vm_group_bin_22697 = frame (4k)
frame_vm_group_bin_22698 = frame (4k)
frame_vm_group_bin_22699 = frame (4k)
frame_vm_group_bin_2270 = frame (4k)
frame_vm_group_bin_22700 = frame (4k)
frame_vm_group_bin_22701 = frame (4k)
frame_vm_group_bin_22702 = frame (4k)
frame_vm_group_bin_22703 = frame (4k)
frame_vm_group_bin_22704 = frame (4k)
frame_vm_group_bin_22705 = frame (4k)
frame_vm_group_bin_22706 = frame (4k)
frame_vm_group_bin_22707 = frame (4k)
frame_vm_group_bin_22708 = frame (4k)
frame_vm_group_bin_22709 = frame (4k)
frame_vm_group_bin_2271 = frame (4k)
frame_vm_group_bin_22710 = frame (4k)
frame_vm_group_bin_22711 = frame (4k)
frame_vm_group_bin_22712 = frame (4k)
frame_vm_group_bin_22713 = frame (4k)
frame_vm_group_bin_22714 = frame (4k)
frame_vm_group_bin_22715 = frame (4k)
frame_vm_group_bin_22716 = frame (4k)
frame_vm_group_bin_22717 = frame (4k)
frame_vm_group_bin_22718 = frame (4k)
frame_vm_group_bin_22719 = frame (4k)
frame_vm_group_bin_2272 = frame (4k)
frame_vm_group_bin_22720 = frame (4k)
frame_vm_group_bin_22721 = frame (4k)
frame_vm_group_bin_22722 = frame (4k)
frame_vm_group_bin_22723 = frame (4k)
frame_vm_group_bin_22724 = frame (4k)
frame_vm_group_bin_22725 = frame (4k)
frame_vm_group_bin_22726 = frame (4k)
frame_vm_group_bin_22727 = frame (4k)
frame_vm_group_bin_22728 = frame (4k)
frame_vm_group_bin_22729 = frame (4k)
frame_vm_group_bin_2273 = frame (4k)
frame_vm_group_bin_22730 = frame (4k)
frame_vm_group_bin_22731 = frame (4k)
frame_vm_group_bin_22732 = frame (4k)
frame_vm_group_bin_22733 = frame (4k)
frame_vm_group_bin_22734 = frame (4k)
frame_vm_group_bin_22735 = frame (4k)
frame_vm_group_bin_22736 = frame (4k)
frame_vm_group_bin_22737 = frame (4k)
frame_vm_group_bin_22738 = frame (4k)
frame_vm_group_bin_22739 = frame (4k)
frame_vm_group_bin_2274 = frame (4k)
frame_vm_group_bin_22740 = frame (4k)
frame_vm_group_bin_22741 = frame (4k)
frame_vm_group_bin_22742 = frame (4k)
frame_vm_group_bin_22743 = frame (4k)
frame_vm_group_bin_22744 = frame (4k)
frame_vm_group_bin_22745 = frame (4k)
frame_vm_group_bin_22746 = frame (4k)
frame_vm_group_bin_22747 = frame (4k)
frame_vm_group_bin_22748 = frame (4k)
frame_vm_group_bin_22749 = frame (4k)
frame_vm_group_bin_2275 = frame (4k)
frame_vm_group_bin_22750 = frame (4k)
frame_vm_group_bin_22751 = frame (4k)
frame_vm_group_bin_22752 = frame (4k)
frame_vm_group_bin_22753 = frame (4k)
frame_vm_group_bin_22754 = frame (4k)
frame_vm_group_bin_22755 = frame (4k)
frame_vm_group_bin_22756 = frame (4k)
frame_vm_group_bin_22757 = frame (4k)
frame_vm_group_bin_22758 = frame (4k)
frame_vm_group_bin_22759 = frame (4k)
frame_vm_group_bin_2276 = frame (4k)
frame_vm_group_bin_22760 = frame (4k)
frame_vm_group_bin_22761 = frame (4k)
frame_vm_group_bin_22762 = frame (4k)
frame_vm_group_bin_22763 = frame (4k)
frame_vm_group_bin_22764 = frame (4k)
frame_vm_group_bin_22765 = frame (4k)
frame_vm_group_bin_22766 = frame (4k)
frame_vm_group_bin_22767 = frame (4k)
frame_vm_group_bin_22768 = frame (4k)
frame_vm_group_bin_22769 = frame (4k)
frame_vm_group_bin_2277 = frame (4k)
frame_vm_group_bin_22770 = frame (4k)
frame_vm_group_bin_22771 = frame (4k)
frame_vm_group_bin_22772 = frame (4k)
frame_vm_group_bin_22773 = frame (4k)
frame_vm_group_bin_22774 = frame (4k)
frame_vm_group_bin_22775 = frame (4k)
frame_vm_group_bin_22776 = frame (4k)
frame_vm_group_bin_22777 = frame (4k)
frame_vm_group_bin_22778 = frame (4k)
frame_vm_group_bin_22779 = frame (4k)
frame_vm_group_bin_2278 = frame (4k)
frame_vm_group_bin_22780 = frame (4k)
frame_vm_group_bin_22781 = frame (4k)
frame_vm_group_bin_22782 = frame (4k)
frame_vm_group_bin_22783 = frame (4k)
frame_vm_group_bin_22784 = frame (4k)
frame_vm_group_bin_22785 = frame (4k)
frame_vm_group_bin_22786 = frame (4k)
frame_vm_group_bin_22787 = frame (4k)
frame_vm_group_bin_22788 = frame (4k)
frame_vm_group_bin_22789 = frame (4k)
frame_vm_group_bin_2279 = frame (4k)
frame_vm_group_bin_22790 = frame (4k)
frame_vm_group_bin_22791 = frame (4k)
frame_vm_group_bin_22792 = frame (4k)
frame_vm_group_bin_22793 = frame (4k)
frame_vm_group_bin_22794 = frame (4k)
frame_vm_group_bin_22795 = frame (4k)
frame_vm_group_bin_22796 = frame (4k)
frame_vm_group_bin_22797 = frame (4k)
frame_vm_group_bin_22798 = frame (4k)
frame_vm_group_bin_22799 = frame (4k)
frame_vm_group_bin_2280 = frame (4k)
frame_vm_group_bin_22800 = frame (4k)
frame_vm_group_bin_22801 = frame (4k)
frame_vm_group_bin_22802 = frame (4k)
frame_vm_group_bin_22803 = frame (4k)
frame_vm_group_bin_22804 = frame (4k)
frame_vm_group_bin_22805 = frame (4k)
frame_vm_group_bin_22806 = frame (4k)
frame_vm_group_bin_22807 = frame (4k)
frame_vm_group_bin_22808 = frame (4k)
frame_vm_group_bin_22809 = frame (4k)
frame_vm_group_bin_2281 = frame (4k)
frame_vm_group_bin_22810 = frame (4k)
frame_vm_group_bin_22811 = frame (4k)
frame_vm_group_bin_22812 = frame (4k)
frame_vm_group_bin_22813 = frame (4k)
frame_vm_group_bin_22814 = frame (4k)
frame_vm_group_bin_22815 = frame (4k)
frame_vm_group_bin_22816 = frame (4k)
frame_vm_group_bin_22817 = frame (4k)
frame_vm_group_bin_22818 = frame (4k)
frame_vm_group_bin_22819 = frame (4k)
frame_vm_group_bin_2282 = frame (4k)
frame_vm_group_bin_22820 = frame (4k)
frame_vm_group_bin_22821 = frame (4k)
frame_vm_group_bin_22822 = frame (4k)
frame_vm_group_bin_22823 = frame (4k)
frame_vm_group_bin_22824 = frame (4k)
frame_vm_group_bin_22825 = frame (4k)
frame_vm_group_bin_22826 = frame (4k)
frame_vm_group_bin_22827 = frame (4k)
frame_vm_group_bin_22828 = frame (4k)
frame_vm_group_bin_22829 = frame (4k)
frame_vm_group_bin_2283 = frame (4k)
frame_vm_group_bin_22830 = frame (4k)
frame_vm_group_bin_22831 = frame (4k)
frame_vm_group_bin_22832 = frame (4k)
frame_vm_group_bin_22833 = frame (4k)
frame_vm_group_bin_22834 = frame (4k)
frame_vm_group_bin_22835 = frame (4k)
frame_vm_group_bin_22836 = frame (4k)
frame_vm_group_bin_22837 = frame (4k)
frame_vm_group_bin_22838 = frame (4k)
frame_vm_group_bin_22839 = frame (4k)
frame_vm_group_bin_2284 = frame (4k)
frame_vm_group_bin_22840 = frame (4k)
frame_vm_group_bin_22841 = frame (4k)
frame_vm_group_bin_22842 = frame (4k)
frame_vm_group_bin_22843 = frame (4k)
frame_vm_group_bin_22844 = frame (4k)
frame_vm_group_bin_22845 = frame (4k)
frame_vm_group_bin_22846 = frame (4k)
frame_vm_group_bin_22847 = frame (4k)
frame_vm_group_bin_22848 = frame (4k)
frame_vm_group_bin_22849 = frame (4k)
frame_vm_group_bin_2285 = frame (4k)
frame_vm_group_bin_22850 = frame (4k)
frame_vm_group_bin_22851 = frame (4k)
frame_vm_group_bin_22852 = frame (4k)
frame_vm_group_bin_22853 = frame (4k)
frame_vm_group_bin_22854 = frame (4k)
frame_vm_group_bin_22855 = frame (4k)
frame_vm_group_bin_22856 = frame (4k)
frame_vm_group_bin_22857 = frame (4k)
frame_vm_group_bin_22858 = frame (4k)
frame_vm_group_bin_22859 = frame (4k)
frame_vm_group_bin_2286 = frame (4k)
frame_vm_group_bin_22860 = frame (4k)
frame_vm_group_bin_22861 = frame (4k)
frame_vm_group_bin_22862 = frame (4k)
frame_vm_group_bin_22863 = frame (4k)
frame_vm_group_bin_22864 = frame (4k)
frame_vm_group_bin_22865 = frame (4k)
frame_vm_group_bin_22866 = frame (4k)
frame_vm_group_bin_22867 = frame (4k)
frame_vm_group_bin_22868 = frame (4k)
frame_vm_group_bin_22869 = frame (4k)
frame_vm_group_bin_2287 = frame (4k)
frame_vm_group_bin_22870 = frame (4k)
frame_vm_group_bin_22871 = frame (4k)
frame_vm_group_bin_22872 = frame (4k)
frame_vm_group_bin_22873 = frame (4k)
frame_vm_group_bin_22874 = frame (4k)
frame_vm_group_bin_22875 = frame (4k)
frame_vm_group_bin_22876 = frame (4k)
frame_vm_group_bin_22877 = frame (4k)
frame_vm_group_bin_22878 = frame (4k)
frame_vm_group_bin_22879 = frame (4k)
frame_vm_group_bin_2288 = frame (4k)
frame_vm_group_bin_22880 = frame (4k)
frame_vm_group_bin_22881 = frame (4k)
frame_vm_group_bin_22882 = frame (4k)
frame_vm_group_bin_22883 = frame (4k)
frame_vm_group_bin_22884 = frame (4k)
frame_vm_group_bin_22885 = frame (4k)
frame_vm_group_bin_22886 = frame (4k)
frame_vm_group_bin_22887 = frame (4k)
frame_vm_group_bin_22888 = frame (4k)
frame_vm_group_bin_22889 = frame (4k)
frame_vm_group_bin_2289 = frame (4k)
frame_vm_group_bin_22890 = frame (4k)
frame_vm_group_bin_22891 = frame (4k)
frame_vm_group_bin_22892 = frame (4k)
frame_vm_group_bin_22893 = frame (4k)
frame_vm_group_bin_22894 = frame (4k)
frame_vm_group_bin_22895 = frame (4k)
frame_vm_group_bin_22896 = frame (4k)
frame_vm_group_bin_22897 = frame (4k)
frame_vm_group_bin_22898 = frame (4k)
frame_vm_group_bin_22899 = frame (4k)
frame_vm_group_bin_2290 = frame (4k)
frame_vm_group_bin_22900 = frame (4k)
frame_vm_group_bin_22901 = frame (4k)
frame_vm_group_bin_22902 = frame (4k)
frame_vm_group_bin_22903 = frame (4k)
frame_vm_group_bin_22904 = frame (4k)
frame_vm_group_bin_22905 = frame (4k)
frame_vm_group_bin_22906 = frame (4k)
frame_vm_group_bin_22907 = frame (4k)
frame_vm_group_bin_22908 = frame (4k)
frame_vm_group_bin_22909 = frame (4k)
frame_vm_group_bin_2291 = frame (4k)
frame_vm_group_bin_22910 = frame (4k)
frame_vm_group_bin_22911 = frame (4k)
frame_vm_group_bin_22912 = frame (4k)
frame_vm_group_bin_22913 = frame (4k)
frame_vm_group_bin_22914 = frame (4k)
frame_vm_group_bin_22915 = frame (4k)
frame_vm_group_bin_22916 = frame (4k)
frame_vm_group_bin_22917 = frame (4k)
frame_vm_group_bin_22918 = frame (4k)
frame_vm_group_bin_22919 = frame (4k)
frame_vm_group_bin_2292 = frame (4k)
frame_vm_group_bin_22920 = frame (4k)
frame_vm_group_bin_22921 = frame (4k)
frame_vm_group_bin_22922 = frame (4k)
frame_vm_group_bin_22923 = frame (4k)
frame_vm_group_bin_22924 = frame (4k)
frame_vm_group_bin_22925 = frame (4k)
frame_vm_group_bin_22926 = frame (4k)
frame_vm_group_bin_22927 = frame (4k)
frame_vm_group_bin_22928 = frame (4k)
frame_vm_group_bin_22929 = frame (4k)
frame_vm_group_bin_2293 = frame (4k)
frame_vm_group_bin_22930 = frame (4k)
frame_vm_group_bin_22931 = frame (4k)
frame_vm_group_bin_22932 = frame (4k)
frame_vm_group_bin_22933 = frame (4k)
frame_vm_group_bin_22934 = frame (4k)
frame_vm_group_bin_22935 = frame (4k)
frame_vm_group_bin_22936 = frame (4k)
frame_vm_group_bin_22937 = frame (4k)
frame_vm_group_bin_22938 = frame (4k)
frame_vm_group_bin_22939 = frame (4k)
frame_vm_group_bin_2294 = frame (4k)
frame_vm_group_bin_22940 = frame (4k)
frame_vm_group_bin_22941 = frame (4k)
frame_vm_group_bin_22942 = frame (4k)
frame_vm_group_bin_22943 = frame (4k)
frame_vm_group_bin_22944 = frame (4k)
frame_vm_group_bin_22945 = frame (4k)
frame_vm_group_bin_22946 = frame (4k)
frame_vm_group_bin_22947 = frame (4k)
frame_vm_group_bin_22948 = frame (4k)
frame_vm_group_bin_22949 = frame (4k)
frame_vm_group_bin_2295 = frame (4k)
frame_vm_group_bin_22950 = frame (4k)
frame_vm_group_bin_22951 = frame (4k)
frame_vm_group_bin_22952 = frame (4k)
frame_vm_group_bin_22953 = frame (4k)
frame_vm_group_bin_22954 = frame (4k)
frame_vm_group_bin_22955 = frame (4k)
frame_vm_group_bin_22956 = frame (4k)
frame_vm_group_bin_22957 = frame (4k)
frame_vm_group_bin_22958 = frame (4k)
frame_vm_group_bin_22959 = frame (4k)
frame_vm_group_bin_2296 = frame (4k)
frame_vm_group_bin_22960 = frame (4k)
frame_vm_group_bin_22961 = frame (4k)
frame_vm_group_bin_22962 = frame (4k)
frame_vm_group_bin_22963 = frame (4k)
frame_vm_group_bin_22964 = frame (4k)
frame_vm_group_bin_22965 = frame (4k)
frame_vm_group_bin_22966 = frame (4k)
frame_vm_group_bin_22967 = frame (4k)
frame_vm_group_bin_22968 = frame (4k)
frame_vm_group_bin_22969 = frame (4k)
frame_vm_group_bin_2297 = frame (4k)
frame_vm_group_bin_22970 = frame (4k)
frame_vm_group_bin_22971 = frame (4k)
frame_vm_group_bin_22972 = frame (4k)
frame_vm_group_bin_22973 = frame (4k)
frame_vm_group_bin_22974 = frame (4k)
frame_vm_group_bin_22975 = frame (4k)
frame_vm_group_bin_22976 = frame (4k)
frame_vm_group_bin_22977 = frame (4k)
frame_vm_group_bin_22978 = frame (4k)
frame_vm_group_bin_22979 = frame (4k)
frame_vm_group_bin_2298 = frame (4k)
frame_vm_group_bin_22980 = frame (4k)
frame_vm_group_bin_22981 = frame (4k)
frame_vm_group_bin_22982 = frame (4k)
frame_vm_group_bin_22983 = frame (4k)
frame_vm_group_bin_22984 = frame (4k)
frame_vm_group_bin_22985 = frame (4k)
frame_vm_group_bin_22986 = frame (4k)
frame_vm_group_bin_22987 = frame (4k)
frame_vm_group_bin_22988 = frame (4k)
frame_vm_group_bin_22989 = frame (4k)
frame_vm_group_bin_2299 = frame (4k)
frame_vm_group_bin_22990 = frame (4k)
frame_vm_group_bin_22991 = frame (4k)
frame_vm_group_bin_22992 = frame (4k)
frame_vm_group_bin_22993 = frame (4k)
frame_vm_group_bin_22994 = frame (4k)
frame_vm_group_bin_22995 = frame (4k)
frame_vm_group_bin_22996 = frame (4k)
frame_vm_group_bin_22997 = frame (4k)
frame_vm_group_bin_22998 = frame (4k)
frame_vm_group_bin_22999 = frame (4k)
frame_vm_group_bin_2300 = frame (4k)
frame_vm_group_bin_23000 = frame (4k)
frame_vm_group_bin_23001 = frame (4k)
frame_vm_group_bin_23002 = frame (4k)
frame_vm_group_bin_23003 = frame (4k)
frame_vm_group_bin_23004 = frame (4k)
frame_vm_group_bin_23005 = frame (4k)
frame_vm_group_bin_23006 = frame (4k)
frame_vm_group_bin_23007 = frame (4k)
frame_vm_group_bin_23008 = frame (4k)
frame_vm_group_bin_23009 = frame (4k)
frame_vm_group_bin_2301 = frame (4k)
frame_vm_group_bin_23010 = frame (4k)
frame_vm_group_bin_23011 = frame (4k)
frame_vm_group_bin_23012 = frame (4k)
frame_vm_group_bin_23013 = frame (4k)
frame_vm_group_bin_23014 = frame (4k)
frame_vm_group_bin_23015 = frame (4k)
frame_vm_group_bin_23016 = frame (4k)
frame_vm_group_bin_23017 = frame (4k)
frame_vm_group_bin_23018 = frame (4k)
frame_vm_group_bin_23019 = frame (4k)
frame_vm_group_bin_2302 = frame (4k)
frame_vm_group_bin_23020 = frame (4k)
frame_vm_group_bin_23021 = frame (4k)
frame_vm_group_bin_23022 = frame (4k)
frame_vm_group_bin_23023 = frame (4k)
frame_vm_group_bin_23024 = frame (4k)
frame_vm_group_bin_23025 = frame (4k)
frame_vm_group_bin_23026 = frame (4k)
frame_vm_group_bin_23027 = frame (4k)
frame_vm_group_bin_23028 = frame (4k)
frame_vm_group_bin_23029 = frame (4k)
frame_vm_group_bin_2303 = frame (4k)
frame_vm_group_bin_23030 = frame (4k)
frame_vm_group_bin_23031 = frame (4k)
frame_vm_group_bin_23032 = frame (4k)
frame_vm_group_bin_23033 = frame (4k)
frame_vm_group_bin_23034 = frame (4k)
frame_vm_group_bin_23035 = frame (4k)
frame_vm_group_bin_23036 = frame (4k)
frame_vm_group_bin_23037 = frame (4k)
frame_vm_group_bin_23038 = frame (4k)
frame_vm_group_bin_23039 = frame (4k)
frame_vm_group_bin_2304 = frame (4k)
frame_vm_group_bin_23040 = frame (4k)
frame_vm_group_bin_23041 = frame (4k)
frame_vm_group_bin_23042 = frame (4k)
frame_vm_group_bin_23043 = frame (4k)
frame_vm_group_bin_23044 = frame (4k)
frame_vm_group_bin_23045 = frame (4k)
frame_vm_group_bin_23046 = frame (4k)
frame_vm_group_bin_23047 = frame (4k)
frame_vm_group_bin_23048 = frame (4k)
frame_vm_group_bin_23049 = frame (4k)
frame_vm_group_bin_2305 = frame (4k)
frame_vm_group_bin_23050 = frame (4k)
frame_vm_group_bin_23051 = frame (4k)
frame_vm_group_bin_23052 = frame (4k)
frame_vm_group_bin_23053 = frame (4k)
frame_vm_group_bin_23054 = frame (4k)
frame_vm_group_bin_23055 = frame (4k)
frame_vm_group_bin_23056 = frame (4k)
frame_vm_group_bin_23057 = frame (4k)
frame_vm_group_bin_23058 = frame (4k)
frame_vm_group_bin_23059 = frame (4k)
frame_vm_group_bin_2306 = frame (4k)
frame_vm_group_bin_23060 = frame (4k)
frame_vm_group_bin_23061 = frame (4k)
frame_vm_group_bin_23062 = frame (4k)
frame_vm_group_bin_23063 = frame (4k)
frame_vm_group_bin_23064 = frame (4k)
frame_vm_group_bin_23065 = frame (4k)
frame_vm_group_bin_23066 = frame (4k)
frame_vm_group_bin_23067 = frame (4k)
frame_vm_group_bin_23068 = frame (4k)
frame_vm_group_bin_23069 = frame (4k)
frame_vm_group_bin_2307 = frame (4k)
frame_vm_group_bin_23070 = frame (4k)
frame_vm_group_bin_23071 = frame (4k)
frame_vm_group_bin_23072 = frame (4k)
frame_vm_group_bin_23073 = frame (4k)
frame_vm_group_bin_23074 = frame (4k)
frame_vm_group_bin_23075 = frame (4k)
frame_vm_group_bin_23076 = frame (4k)
frame_vm_group_bin_23077 = frame (4k)
frame_vm_group_bin_23078 = frame (4k)
frame_vm_group_bin_23079 = frame (4k)
frame_vm_group_bin_2308 = frame (4k)
frame_vm_group_bin_23080 = frame (4k)
frame_vm_group_bin_23081 = frame (4k)
frame_vm_group_bin_23082 = frame (4k)
frame_vm_group_bin_23083 = frame (4k)
frame_vm_group_bin_23084 = frame (4k)
frame_vm_group_bin_23085 = frame (4k)
frame_vm_group_bin_23086 = frame (4k)
frame_vm_group_bin_23087 = frame (4k)
frame_vm_group_bin_23088 = frame (4k)
frame_vm_group_bin_23089 = frame (4k)
frame_vm_group_bin_2309 = frame (4k)
frame_vm_group_bin_23090 = frame (4k)
frame_vm_group_bin_23091 = frame (4k)
frame_vm_group_bin_23092 = frame (4k)
frame_vm_group_bin_23093 = frame (4k)
frame_vm_group_bin_23094 = frame (4k)
frame_vm_group_bin_23095 = frame (4k)
frame_vm_group_bin_23096 = frame (4k)
frame_vm_group_bin_23097 = frame (4k)
frame_vm_group_bin_23098 = frame (4k)
frame_vm_group_bin_23099 = frame (4k)
frame_vm_group_bin_2310 = frame (4k)
frame_vm_group_bin_23100 = frame (4k)
frame_vm_group_bin_23101 = frame (4k)
frame_vm_group_bin_23102 = frame (4k)
frame_vm_group_bin_23103 = frame (4k)
frame_vm_group_bin_23104 = frame (4k)
frame_vm_group_bin_23105 = frame (4k)
frame_vm_group_bin_23106 = frame (4k)
frame_vm_group_bin_23107 = frame (4k)
frame_vm_group_bin_23108 = frame (4k)
frame_vm_group_bin_23109 = frame (4k)
frame_vm_group_bin_2311 = frame (4k)
frame_vm_group_bin_23110 = frame (4k)
frame_vm_group_bin_23111 = frame (4k)
frame_vm_group_bin_23112 = frame (4k)
frame_vm_group_bin_23113 = frame (4k)
frame_vm_group_bin_23114 = frame (4k)
frame_vm_group_bin_23115 = frame (4k)
frame_vm_group_bin_23116 = frame (4k)
frame_vm_group_bin_23117 = frame (4k)
frame_vm_group_bin_23118 = frame (4k)
frame_vm_group_bin_23119 = frame (4k)
frame_vm_group_bin_2312 = frame (4k)
frame_vm_group_bin_23120 = frame (4k)
frame_vm_group_bin_23121 = frame (4k)
frame_vm_group_bin_23122 = frame (4k)
frame_vm_group_bin_23123 = frame (4k)
frame_vm_group_bin_23124 = frame (4k)
frame_vm_group_bin_23125 = frame (4k)
frame_vm_group_bin_23126 = frame (4k)
frame_vm_group_bin_23127 = frame (4k)
frame_vm_group_bin_23128 = frame (4k)
frame_vm_group_bin_23129 = frame (4k)
frame_vm_group_bin_2313 = frame (4k)
frame_vm_group_bin_23130 = frame (4k)
frame_vm_group_bin_23131 = frame (4k)
frame_vm_group_bin_23132 = frame (4k)
frame_vm_group_bin_23133 = frame (4k)
frame_vm_group_bin_23134 = frame (4k)
frame_vm_group_bin_23135 = frame (4k)
frame_vm_group_bin_23136 = frame (4k)
frame_vm_group_bin_23137 = frame (4k)
frame_vm_group_bin_23138 = frame (4k)
frame_vm_group_bin_23139 = frame (4k)
frame_vm_group_bin_2314 = frame (4k)
frame_vm_group_bin_23140 = frame (4k)
frame_vm_group_bin_23141 = frame (4k)
frame_vm_group_bin_23142 = frame (4k)
frame_vm_group_bin_23143 = frame (4k)
frame_vm_group_bin_23144 = frame (4k)
frame_vm_group_bin_23145 = frame (4k)
frame_vm_group_bin_23146 = frame (4k)
frame_vm_group_bin_23147 = frame (4k)
frame_vm_group_bin_23148 = frame (4k)
frame_vm_group_bin_23149 = frame (4k)
frame_vm_group_bin_2315 = frame (4k)
frame_vm_group_bin_23150 = frame (4k)
frame_vm_group_bin_23151 = frame (4k)
frame_vm_group_bin_23152 = frame (4k)
frame_vm_group_bin_23153 = frame (4k)
frame_vm_group_bin_23154 = frame (4k)
frame_vm_group_bin_23155 = frame (4k)
frame_vm_group_bin_23156 = frame (4k)
frame_vm_group_bin_23157 = frame (4k)
frame_vm_group_bin_23158 = frame (4k)
frame_vm_group_bin_23159 = frame (4k)
frame_vm_group_bin_2316 = frame (4k)
frame_vm_group_bin_23160 = frame (4k)
frame_vm_group_bin_23161 = frame (4k)
frame_vm_group_bin_23162 = frame (4k)
frame_vm_group_bin_23163 = frame (4k)
frame_vm_group_bin_23164 = frame (4k)
frame_vm_group_bin_23165 = frame (4k)
frame_vm_group_bin_23166 = frame (4k)
frame_vm_group_bin_23167 = frame (4k)
frame_vm_group_bin_23168 = frame (4k)
frame_vm_group_bin_23169 = frame (4k)
frame_vm_group_bin_2317 = frame (4k)
frame_vm_group_bin_23170 = frame (4k)
frame_vm_group_bin_23171 = frame (4k)
frame_vm_group_bin_23172 = frame (4k)
frame_vm_group_bin_23173 = frame (4k)
frame_vm_group_bin_23174 = frame (4k)
frame_vm_group_bin_23175 = frame (4k)
frame_vm_group_bin_23176 = frame (4k)
frame_vm_group_bin_23177 = frame (4k)
frame_vm_group_bin_23178 = frame (4k)
frame_vm_group_bin_23179 = frame (4k)
frame_vm_group_bin_2318 = frame (4k)
frame_vm_group_bin_23180 = frame (4k)
frame_vm_group_bin_23181 = frame (4k)
frame_vm_group_bin_23182 = frame (4k)
frame_vm_group_bin_23183 = frame (4k)
frame_vm_group_bin_23184 = frame (4k)
frame_vm_group_bin_23185 = frame (4k)
frame_vm_group_bin_23186 = frame (4k)
frame_vm_group_bin_23187 = frame (4k)
frame_vm_group_bin_23188 = frame (4k)
frame_vm_group_bin_23189 = frame (4k)
frame_vm_group_bin_2319 = frame (4k)
frame_vm_group_bin_23190 = frame (4k)
frame_vm_group_bin_23191 = frame (4k)
frame_vm_group_bin_23192 = frame (4k)
frame_vm_group_bin_23193 = frame (4k)
frame_vm_group_bin_23195 = frame (4k)
frame_vm_group_bin_23196 = frame (4k)
frame_vm_group_bin_23197 = frame (4k)
frame_vm_group_bin_23198 = frame (4k)
frame_vm_group_bin_23199 = frame (4k)
frame_vm_group_bin_2320 = frame (4k)
frame_vm_group_bin_23200 = frame (4k)
frame_vm_group_bin_23201 = frame (4k)
frame_vm_group_bin_23202 = frame (4k)
frame_vm_group_bin_23203 = frame (4k)
frame_vm_group_bin_23204 = frame (4k)
frame_vm_group_bin_23205 = frame (4k)
frame_vm_group_bin_23206 = frame (4k)
frame_vm_group_bin_23207 = frame (4k)
frame_vm_group_bin_23208 = frame (4k)
frame_vm_group_bin_23209 = frame (4k)
frame_vm_group_bin_2321 = frame (4k)
frame_vm_group_bin_23210 = frame (4k)
frame_vm_group_bin_23211 = frame (4k)
frame_vm_group_bin_23212 = frame (4k)
frame_vm_group_bin_23213 = frame (4k)
frame_vm_group_bin_23214 = frame (4k)
frame_vm_group_bin_23215 = frame (4k)
frame_vm_group_bin_23216 = frame (4k)
frame_vm_group_bin_23217 = frame (4k)
frame_vm_group_bin_23218 = frame (4k)
frame_vm_group_bin_23219 = frame (4k)
frame_vm_group_bin_2322 = frame (4k)
frame_vm_group_bin_23220 = frame (4k)
frame_vm_group_bin_23221 = frame (4k)
frame_vm_group_bin_23222 = frame (4k)
frame_vm_group_bin_23223 = frame (4k)
frame_vm_group_bin_23224 = frame (4k)
frame_vm_group_bin_23225 = frame (4k)
frame_vm_group_bin_23226 = frame (4k)
frame_vm_group_bin_23227 = frame (4k)
frame_vm_group_bin_23228 = frame (4k)
frame_vm_group_bin_23229 = frame (4k)
frame_vm_group_bin_2323 = frame (4k)
frame_vm_group_bin_23230 = frame (4k)
frame_vm_group_bin_23231 = frame (4k)
frame_vm_group_bin_23232 = frame (4k)
frame_vm_group_bin_23233 = frame (4k)
frame_vm_group_bin_23234 = frame (4k)
frame_vm_group_bin_23235 = frame (4k)
frame_vm_group_bin_23236 = frame (4k)
frame_vm_group_bin_23237 = frame (4k)
frame_vm_group_bin_23238 = frame (4k)
frame_vm_group_bin_23239 = frame (4k)
frame_vm_group_bin_2324 = frame (4k)
frame_vm_group_bin_23240 = frame (4k)
frame_vm_group_bin_23241 = frame (4k)
frame_vm_group_bin_23242 = frame (4k)
frame_vm_group_bin_23243 = frame (4k)
frame_vm_group_bin_23244 = frame (4k)
frame_vm_group_bin_23245 = frame (4k)
frame_vm_group_bin_23246 = frame (4k)
frame_vm_group_bin_23247 = frame (4k)
frame_vm_group_bin_23248 = frame (4k)
frame_vm_group_bin_23249 = frame (4k)
frame_vm_group_bin_2325 = frame (4k)
frame_vm_group_bin_23250 = frame (4k)
frame_vm_group_bin_23251 = frame (4k)
frame_vm_group_bin_23252 = frame (4k)
frame_vm_group_bin_23253 = frame (4k)
frame_vm_group_bin_23254 = frame (4k)
frame_vm_group_bin_23255 = frame (4k)
frame_vm_group_bin_2326 = frame (4k)
frame_vm_group_bin_2327 = frame (4k)
frame_vm_group_bin_2328 = frame (4k)
frame_vm_group_bin_2329 = frame (4k)
frame_vm_group_bin_2330 = frame (4k)
frame_vm_group_bin_2331 = frame (4k)
frame_vm_group_bin_2332 = frame (4k)
frame_vm_group_bin_2333 = frame (4k)
frame_vm_group_bin_2334 = frame (4k)
frame_vm_group_bin_2335 = frame (4k)
frame_vm_group_bin_2336 = frame (4k)
frame_vm_group_bin_2337 = frame (4k)
frame_vm_group_bin_2338 = frame (4k)
frame_vm_group_bin_2339 = frame (4k)
frame_vm_group_bin_2340 = frame (4k)
frame_vm_group_bin_2341 = frame (4k)
frame_vm_group_bin_2342 = frame (4k)
frame_vm_group_bin_2343 = frame (4k)
frame_vm_group_bin_2344 = frame (4k)
frame_vm_group_bin_2345 = frame (4k)
frame_vm_group_bin_2346 = frame (4k)
frame_vm_group_bin_2347 = frame (4k)
frame_vm_group_bin_2348 = frame (4k)
frame_vm_group_bin_2349 = frame (4k)
frame_vm_group_bin_2350 = frame (4k)
frame_vm_group_bin_2351 = frame (4k)
frame_vm_group_bin_2352 = frame (4k)
frame_vm_group_bin_2353 = frame (4k)
frame_vm_group_bin_2354 = frame (4k)
frame_vm_group_bin_2355 = frame (4k)
frame_vm_group_bin_2356 = frame (4k)
frame_vm_group_bin_2357 = frame (4k)
frame_vm_group_bin_2358 = frame (4k)
frame_vm_group_bin_2359 = frame (4k)
frame_vm_group_bin_2360 = frame (4k)
frame_vm_group_bin_2361 = frame (4k)
frame_vm_group_bin_2362 = frame (4k)
frame_vm_group_bin_2363 = frame (4k)
frame_vm_group_bin_2364 = frame (4k)
frame_vm_group_bin_2365 = frame (4k)
frame_vm_group_bin_2366 = frame (4k)
frame_vm_group_bin_2367 = frame (4k)
frame_vm_group_bin_2368 = frame (4k)
frame_vm_group_bin_2369 = frame (4k)
frame_vm_group_bin_2370 = frame (4k)
frame_vm_group_bin_2371 = frame (4k)
frame_vm_group_bin_2372 = frame (4k)
frame_vm_group_bin_2373 = frame (4k)
frame_vm_group_bin_2374 = frame (4k)
frame_vm_group_bin_2375 = frame (4k)
frame_vm_group_bin_2376 = frame (4k)
frame_vm_group_bin_2377 = frame (4k)
frame_vm_group_bin_2378 = frame (4k)
frame_vm_group_bin_2379 = frame (4k)
frame_vm_group_bin_2380 = frame (4k)
frame_vm_group_bin_2381 = frame (4k)
frame_vm_group_bin_2382 = frame (4k)
frame_vm_group_bin_2383 = frame (4k)
frame_vm_group_bin_2384 = frame (4k)
frame_vm_group_bin_2385 = frame (4k)
frame_vm_group_bin_2386 = frame (4k)
frame_vm_group_bin_2387 = frame (4k)
frame_vm_group_bin_2388 = frame (4k)
frame_vm_group_bin_2389 = frame (4k)
frame_vm_group_bin_2390 = frame (4k)
frame_vm_group_bin_2391 = frame (4k)
frame_vm_group_bin_2392 = frame (4k)
frame_vm_group_bin_2393 = frame (4k)
frame_vm_group_bin_2394 = frame (4k)
frame_vm_group_bin_2395 = frame (4k)
frame_vm_group_bin_2396 = frame (4k)
frame_vm_group_bin_2397 = frame (4k)
frame_vm_group_bin_2398 = frame (4k)
frame_vm_group_bin_2399 = frame (4k)
frame_vm_group_bin_2400 = frame (4k)
frame_vm_group_bin_2401 = frame (4k)
frame_vm_group_bin_2402 = frame (4k)
frame_vm_group_bin_2403 = frame (4k)
frame_vm_group_bin_2404 = frame (4k)
frame_vm_group_bin_2405 = frame (4k)
frame_vm_group_bin_2406 = frame (4k)
frame_vm_group_bin_2407 = frame (4k)
frame_vm_group_bin_2408 = frame (4k)
frame_vm_group_bin_2409 = frame (4k)
frame_vm_group_bin_2410 = frame (4k)
frame_vm_group_bin_2411 = frame (4k)
frame_vm_group_bin_2412 = frame (4k)
frame_vm_group_bin_2413 = frame (4k)
frame_vm_group_bin_2414 = frame (4k)
frame_vm_group_bin_2415 = frame (4k)
frame_vm_group_bin_2416 = frame (4k)
frame_vm_group_bin_2417 = frame (4k)
frame_vm_group_bin_2418 = frame (4k)
frame_vm_group_bin_2419 = frame (4k)
frame_vm_group_bin_2420 = frame (4k)
frame_vm_group_bin_2421 = frame (4k)
frame_vm_group_bin_2422 = frame (4k)
frame_vm_group_bin_2423 = frame (4k)
frame_vm_group_bin_2424 = frame (4k)
frame_vm_group_bin_2425 = frame (4k)
frame_vm_group_bin_2426 = frame (4k)
frame_vm_group_bin_2427 = frame (4k)
frame_vm_group_bin_2428 = frame (4k)
frame_vm_group_bin_2429 = frame (4k)
frame_vm_group_bin_2430 = frame (4k)
frame_vm_group_bin_2431 = frame (4k)
frame_vm_group_bin_2432 = frame (4k)
frame_vm_group_bin_2433 = frame (4k)
frame_vm_group_bin_2434 = frame (4k)
frame_vm_group_bin_2435 = frame (4k)
frame_vm_group_bin_2436 = frame (4k)
frame_vm_group_bin_2437 = frame (4k)
frame_vm_group_bin_2438 = frame (4k)
frame_vm_group_bin_2439 = frame (4k)
frame_vm_group_bin_2440 = frame (4k)
frame_vm_group_bin_2441 = frame (4k)
frame_vm_group_bin_2442 = frame (4k)
frame_vm_group_bin_2443 = frame (4k)
frame_vm_group_bin_2444 = frame (4k)
frame_vm_group_bin_2445 = frame (4k)
frame_vm_group_bin_2446 = frame (4k)
frame_vm_group_bin_2447 = frame (4k)
frame_vm_group_bin_2448 = frame (4k)
frame_vm_group_bin_2449 = frame (4k)
frame_vm_group_bin_2450 = frame (4k)
frame_vm_group_bin_2451 = frame (4k)
frame_vm_group_bin_2452 = frame (4k)
frame_vm_group_bin_2453 = frame (4k)
frame_vm_group_bin_2454 = frame (4k)
frame_vm_group_bin_2455 = frame (4k)
frame_vm_group_bin_2456 = frame (4k)
frame_vm_group_bin_2457 = frame (4k)
frame_vm_group_bin_2458 = frame (4k)
frame_vm_group_bin_2459 = frame (4k)
frame_vm_group_bin_2460 = frame (4k)
frame_vm_group_bin_2461 = frame (4k)
frame_vm_group_bin_2462 = frame (4k)
frame_vm_group_bin_2463 = frame (4k)
frame_vm_group_bin_2464 = frame (4k)
frame_vm_group_bin_2465 = frame (4k)
frame_vm_group_bin_2466 = frame (4k)
frame_vm_group_bin_2467 = frame (4k)
frame_vm_group_bin_2468 = frame (4k)
frame_vm_group_bin_2469 = frame (4k)
frame_vm_group_bin_2470 = frame (4k)
frame_vm_group_bin_2471 = frame (4k)
frame_vm_group_bin_2472 = frame (4k)
frame_vm_group_bin_2473 = frame (4k)
frame_vm_group_bin_2474 = frame (4k)
frame_vm_group_bin_2475 = frame (4k)
frame_vm_group_bin_2476 = frame (4k)
frame_vm_group_bin_2477 = frame (4k)
frame_vm_group_bin_2478 = frame (4k)
frame_vm_group_bin_2479 = frame (4k)
frame_vm_group_bin_2480 = frame (4k)
frame_vm_group_bin_2481 = frame (4k)
frame_vm_group_bin_2482 = frame (4k)
frame_vm_group_bin_2483 = frame (4k)
frame_vm_group_bin_2484 = frame (4k)
frame_vm_group_bin_2485 = frame (4k)
frame_vm_group_bin_2486 = frame (4k)
frame_vm_group_bin_2487 = frame (4k)
frame_vm_group_bin_2488 = frame (4k)
frame_vm_group_bin_2489 = frame (4k)
frame_vm_group_bin_2490 = frame (4k)
frame_vm_group_bin_2491 = frame (4k)
frame_vm_group_bin_2492 = frame (4k)
frame_vm_group_bin_2493 = frame (4k)
frame_vm_group_bin_2494 = frame (4k)
frame_vm_group_bin_2495 = frame (4k)
frame_vm_group_bin_2496 = frame (4k)
frame_vm_group_bin_2497 = frame (4k)
frame_vm_group_bin_2498 = frame (4k)
frame_vm_group_bin_2499 = frame (4k)
frame_vm_group_bin_2500 = frame (4k)
frame_vm_group_bin_2501 = frame (4k)
frame_vm_group_bin_2502 = frame (4k)
frame_vm_group_bin_2503 = frame (4k)
frame_vm_group_bin_2504 = frame (4k)
frame_vm_group_bin_2505 = frame (4k)
frame_vm_group_bin_2506 = frame (4k)
frame_vm_group_bin_2507 = frame (4k)
frame_vm_group_bin_2508 = frame (4k)
frame_vm_group_bin_2509 = frame (4k)
frame_vm_group_bin_2510 = frame (4k)
frame_vm_group_bin_2511 = frame (4k)
frame_vm_group_bin_2512 = frame (4k)
frame_vm_group_bin_2513 = frame (4k)
frame_vm_group_bin_2514 = frame (4k)
frame_vm_group_bin_2515 = frame (4k)
frame_vm_group_bin_2516 = frame (4k)
frame_vm_group_bin_2517 = frame (4k)
frame_vm_group_bin_2518 = frame (4k)
frame_vm_group_bin_2519 = frame (4k)
frame_vm_group_bin_2520 = frame (4k)
frame_vm_group_bin_2521 = frame (4k)
frame_vm_group_bin_2522 = frame (4k)
frame_vm_group_bin_2523 = frame (4k)
frame_vm_group_bin_2524 = frame (4k)
frame_vm_group_bin_2525 = frame (4k)
frame_vm_group_bin_2526 = frame (4k)
frame_vm_group_bin_2527 = frame (4k)
frame_vm_group_bin_2528 = frame (4k)
frame_vm_group_bin_2529 = frame (4k)
frame_vm_group_bin_2530 = frame (4k)
frame_vm_group_bin_2531 = frame (4k)
frame_vm_group_bin_2532 = frame (4k)
frame_vm_group_bin_2533 = frame (4k)
frame_vm_group_bin_2534 = frame (4k)
frame_vm_group_bin_2535 = frame (4k)
frame_vm_group_bin_2536 = frame (4k)
frame_vm_group_bin_2537 = frame (4k)
frame_vm_group_bin_2538 = frame (4k)
frame_vm_group_bin_2539 = frame (4k)
frame_vm_group_bin_2540 = frame (4k)
frame_vm_group_bin_2541 = frame (4k)
frame_vm_group_bin_2542 = frame (4k)
frame_vm_group_bin_2543 = frame (4k)
frame_vm_group_bin_2544 = frame (4k)
frame_vm_group_bin_2545 = frame (4k)
frame_vm_group_bin_2546 = frame (4k)
frame_vm_group_bin_2547 = frame (4k)
frame_vm_group_bin_2548 = frame (4k)
frame_vm_group_bin_2549 = frame (4k)
frame_vm_group_bin_2550 = frame (4k)
frame_vm_group_bin_2551 = frame (4k)
frame_vm_group_bin_2552 = frame (4k)
frame_vm_group_bin_2553 = frame (4k)
frame_vm_group_bin_2554 = frame (4k)
frame_vm_group_bin_2555 = frame (4k)
frame_vm_group_bin_2556 = frame (4k)
frame_vm_group_bin_2557 = frame (4k)
frame_vm_group_bin_2558 = frame (4k)
frame_vm_group_bin_2559 = frame (4k)
frame_vm_group_bin_2560 = frame (4k)
frame_vm_group_bin_2561 = frame (4k)
frame_vm_group_bin_2562 = frame (4k)
frame_vm_group_bin_2563 = frame (4k)
frame_vm_group_bin_2564 = frame (4k)
frame_vm_group_bin_2565 = frame (4k)
frame_vm_group_bin_2566 = frame (4k)
frame_vm_group_bin_2567 = frame (4k)
frame_vm_group_bin_2568 = frame (4k)
frame_vm_group_bin_2569 = frame (4k)
frame_vm_group_bin_2570 = frame (4k)
frame_vm_group_bin_2571 = frame (4k)
frame_vm_group_bin_2572 = frame (4k)
frame_vm_group_bin_2573 = frame (4k)
frame_vm_group_bin_2574 = frame (4k)
frame_vm_group_bin_2575 = frame (4k)
frame_vm_group_bin_2576 = frame (4k)
frame_vm_group_bin_2577 = frame (4k)
frame_vm_group_bin_2578 = frame (4k)
frame_vm_group_bin_2579 = frame (4k)
frame_vm_group_bin_2580 = frame (4k)
frame_vm_group_bin_2581 = frame (4k)
frame_vm_group_bin_2582 = frame (4k)
frame_vm_group_bin_2583 = frame (4k)
frame_vm_group_bin_2584 = frame (4k)
frame_vm_group_bin_2585 = frame (4k)
frame_vm_group_bin_2586 = frame (4k)
frame_vm_group_bin_2587 = frame (4k)
frame_vm_group_bin_2588 = frame (4k)
frame_vm_group_bin_2589 = frame (4k)
frame_vm_group_bin_2590 = frame (4k)
frame_vm_group_bin_2591 = frame (4k)
frame_vm_group_bin_2592 = frame (4k)
frame_vm_group_bin_2593 = frame (4k)
frame_vm_group_bin_2594 = frame (4k)
frame_vm_group_bin_2595 = frame (4k)
frame_vm_group_bin_2596 = frame (4k)
frame_vm_group_bin_2597 = frame (4k)
frame_vm_group_bin_2598 = frame (4k)
frame_vm_group_bin_2599 = frame (4k)
frame_vm_group_bin_2600 = frame (4k)
frame_vm_group_bin_2601 = frame (4k)
frame_vm_group_bin_2602 = frame (4k)
frame_vm_group_bin_2603 = frame (4k)
frame_vm_group_bin_2604 = frame (4k)
frame_vm_group_bin_2605 = frame (4k)
frame_vm_group_bin_2606 = frame (4k)
frame_vm_group_bin_2607 = frame (4k)
frame_vm_group_bin_2608 = frame (4k)
frame_vm_group_bin_2609 = frame (4k)
frame_vm_group_bin_2610 = frame (4k)
frame_vm_group_bin_2611 = frame (4k)
frame_vm_group_bin_2612 = frame (4k)
frame_vm_group_bin_2613 = frame (4k)
frame_vm_group_bin_2614 = frame (4k)
frame_vm_group_bin_2615 = frame (4k)
frame_vm_group_bin_2616 = frame (4k)
frame_vm_group_bin_2617 = frame (4k)
frame_vm_group_bin_2618 = frame (4k)
frame_vm_group_bin_2619 = frame (4k)
frame_vm_group_bin_2620 = frame (4k)
frame_vm_group_bin_2621 = frame (4k)
frame_vm_group_bin_2622 = frame (4k)
frame_vm_group_bin_2623 = frame (4k)
frame_vm_group_bin_2624 = frame (4k)
frame_vm_group_bin_2625 = frame (4k)
frame_vm_group_bin_2626 = frame (4k)
frame_vm_group_bin_2627 = frame (4k)
frame_vm_group_bin_2628 = frame (4k)
frame_vm_group_bin_2629 = frame (4k)
frame_vm_group_bin_2630 = frame (4k)
frame_vm_group_bin_2631 = frame (4k)
frame_vm_group_bin_2632 = frame (4k)
frame_vm_group_bin_2633 = frame (4k)
frame_vm_group_bin_2634 = frame (4k)
frame_vm_group_bin_2635 = frame (4k)
frame_vm_group_bin_2636 = frame (4k)
frame_vm_group_bin_2637 = frame (4k)
frame_vm_group_bin_2638 = frame (4k)
frame_vm_group_bin_2639 = frame (4k)
frame_vm_group_bin_2640 = frame (4k)
frame_vm_group_bin_2641 = frame (4k)
frame_vm_group_bin_2642 = frame (4k)
frame_vm_group_bin_2643 = frame (4k)
frame_vm_group_bin_2644 = frame (4k)
frame_vm_group_bin_2645 = frame (4k)
frame_vm_group_bin_2646 = frame (4k)
frame_vm_group_bin_2647 = frame (4k)
frame_vm_group_bin_2648 = frame (4k)
frame_vm_group_bin_2649 = frame (4k)
frame_vm_group_bin_2650 = frame (4k)
frame_vm_group_bin_2651 = frame (4k)
frame_vm_group_bin_2652 = frame (4k)
frame_vm_group_bin_2653 = frame (4k)
frame_vm_group_bin_2654 = frame (4k)
frame_vm_group_bin_2655 = frame (4k)
frame_vm_group_bin_2656 = frame (4k)
frame_vm_group_bin_2657 = frame (4k)
frame_vm_group_bin_2658 = frame (4k)
frame_vm_group_bin_2659 = frame (4k)
frame_vm_group_bin_2660 = frame (4k)
frame_vm_group_bin_2661 = frame (4k)
frame_vm_group_bin_2662 = frame (4k)
frame_vm_group_bin_2663 = frame (4k)
frame_vm_group_bin_2664 = frame (4k)
frame_vm_group_bin_2665 = frame (4k)
frame_vm_group_bin_2666 = frame (4k)
frame_vm_group_bin_2667 = frame (4k)
frame_vm_group_bin_2668 = frame (4k)
frame_vm_group_bin_2669 = frame (4k)
frame_vm_group_bin_2670 = frame (4k)
frame_vm_group_bin_2671 = frame (4k)
frame_vm_group_bin_2672 = frame (4k)
frame_vm_group_bin_2673 = frame (4k)
frame_vm_group_bin_2674 = frame (4k)
frame_vm_group_bin_2675 = frame (4k)
frame_vm_group_bin_2676 = frame (4k)
frame_vm_group_bin_2677 = frame (4k)
frame_vm_group_bin_2678 = frame (4k)
frame_vm_group_bin_2679 = frame (4k)
frame_vm_group_bin_2680 = frame (4k)
frame_vm_group_bin_2681 = frame (4k)
frame_vm_group_bin_2682 = frame (4k)
frame_vm_group_bin_2683 = frame (4k)
frame_vm_group_bin_2684 = frame (4k)
frame_vm_group_bin_2685 = frame (4k)
frame_vm_group_bin_2686 = frame (4k)
frame_vm_group_bin_2687 = frame (4k)
frame_vm_group_bin_2688 = frame (4k)
frame_vm_group_bin_2689 = frame (4k)
frame_vm_group_bin_2690 = frame (4k)
frame_vm_group_bin_2691 = frame (4k)
frame_vm_group_bin_2692 = frame (4k)
frame_vm_group_bin_2693 = frame (4k)
frame_vm_group_bin_2694 = frame (4k)
frame_vm_group_bin_2695 = frame (4k)
frame_vm_group_bin_2696 = frame (4k)
frame_vm_group_bin_2697 = frame (4k)
frame_vm_group_bin_2698 = frame (4k)
frame_vm_group_bin_2699 = frame (4k)
frame_vm_group_bin_2700 = frame (4k)
frame_vm_group_bin_2701 = frame (4k)
frame_vm_group_bin_2702 = frame (4k)
frame_vm_group_bin_2703 = frame (4k)
frame_vm_group_bin_2704 = frame (4k)
frame_vm_group_bin_2705 = frame (4k)
frame_vm_group_bin_2706 = frame (4k)
frame_vm_group_bin_2707 = frame (4k)
frame_vm_group_bin_2708 = frame (4k)
frame_vm_group_bin_2709 = frame (4k)
frame_vm_group_bin_2710 = frame (4k)
frame_vm_group_bin_2711 = frame (4k)
frame_vm_group_bin_2712 = frame (4k)
frame_vm_group_bin_2713 = frame (4k)
frame_vm_group_bin_2714 = frame (4k)
frame_vm_group_bin_2715 = frame (4k)
frame_vm_group_bin_2716 = frame (4k)
frame_vm_group_bin_2717 = frame (4k)
frame_vm_group_bin_2718 = frame (4k)
frame_vm_group_bin_2719 = frame (4k)
frame_vm_group_bin_2720 = frame (4k)
frame_vm_group_bin_2721 = frame (4k)
frame_vm_group_bin_2722 = frame (4k)
frame_vm_group_bin_2723 = frame (4k)
frame_vm_group_bin_2724 = frame (4k)
frame_vm_group_bin_2725 = frame (4k)
frame_vm_group_bin_2726 = frame (4k)
frame_vm_group_bin_2727 = frame (4k)
frame_vm_group_bin_2728 = frame (4k)
frame_vm_group_bin_2729 = frame (4k)
frame_vm_group_bin_2730 = frame (4k)
frame_vm_group_bin_2731 = frame (4k)
frame_vm_group_bin_2732 = frame (4k)
frame_vm_group_bin_2733 = frame (4k)
frame_vm_group_bin_2734 = frame (4k)
frame_vm_group_bin_2735 = frame (4k)
frame_vm_group_bin_2736 = frame (4k)
frame_vm_group_bin_2737 = frame (4k)
frame_vm_group_bin_2738 = frame (4k)
frame_vm_group_bin_2739 = frame (4k)
frame_vm_group_bin_2740 = frame (4k)
frame_vm_group_bin_2741 = frame (4k)
frame_vm_group_bin_2742 = frame (4k)
frame_vm_group_bin_2743 = frame (4k)
frame_vm_group_bin_2744 = frame (4k)
frame_vm_group_bin_2745 = frame (4k)
frame_vm_group_bin_2746 = frame (4k)
frame_vm_group_bin_2747 = frame (4k)
frame_vm_group_bin_2748 = frame (4k)
frame_vm_group_bin_2749 = frame (4k)
frame_vm_group_bin_2750 = frame (4k)
frame_vm_group_bin_2751 = frame (4k)
frame_vm_group_bin_2752 = frame (4k)
frame_vm_group_bin_2753 = frame (4k)
frame_vm_group_bin_2754 = frame (4k)
frame_vm_group_bin_2755 = frame (4k)
frame_vm_group_bin_2756 = frame (4k)
frame_vm_group_bin_2757 = frame (4k)
frame_vm_group_bin_2758 = frame (4k)
frame_vm_group_bin_2759 = frame (4k)
frame_vm_group_bin_2760 = frame (4k)
frame_vm_group_bin_2761 = frame (4k)
frame_vm_group_bin_2762 = frame (4k)
frame_vm_group_bin_2763 = frame (4k)
frame_vm_group_bin_2764 = frame (4k)
frame_vm_group_bin_2765 = frame (4k)
frame_vm_group_bin_2766 = frame (4k)
frame_vm_group_bin_2767 = frame (4k)
frame_vm_group_bin_2768 = frame (4k)
frame_vm_group_bin_2769 = frame (4k)
frame_vm_group_bin_2770 = frame (4k)
frame_vm_group_bin_2771 = frame (4k)
frame_vm_group_bin_2772 = frame (4k)
frame_vm_group_bin_2773 = frame (4k)
frame_vm_group_bin_2774 = frame (4k)
frame_vm_group_bin_2775 = frame (4k)
frame_vm_group_bin_2776 = frame (4k)
frame_vm_group_bin_2777 = frame (4k)
frame_vm_group_bin_2778 = frame (4k)
frame_vm_group_bin_2779 = frame (4k)
frame_vm_group_bin_2780 = frame (4k)
frame_vm_group_bin_2781 = frame (4k)
frame_vm_group_bin_2782 = frame (4k)
frame_vm_group_bin_2783 = frame (4k)
frame_vm_group_bin_2784 = frame (4k)
frame_vm_group_bin_2785 = frame (4k)
frame_vm_group_bin_2786 = frame (4k)
frame_vm_group_bin_2787 = frame (4k)
frame_vm_group_bin_2788 = frame (4k)
frame_vm_group_bin_2789 = frame (4k)
frame_vm_group_bin_2790 = frame (4k)
frame_vm_group_bin_2791 = frame (4k)
frame_vm_group_bin_2792 = frame (4k)
frame_vm_group_bin_2793 = frame (4k)
frame_vm_group_bin_2794 = frame (4k)
frame_vm_group_bin_2795 = frame (4k)
frame_vm_group_bin_2796 = frame (4k)
frame_vm_group_bin_2797 = frame (4k)
frame_vm_group_bin_2798 = frame (4k)
frame_vm_group_bin_2799 = frame (4k)
frame_vm_group_bin_2800 = frame (4k)
frame_vm_group_bin_2801 = frame (4k)
frame_vm_group_bin_2802 = frame (4k)
frame_vm_group_bin_2803 = frame (4k)
frame_vm_group_bin_2804 = frame (4k)
frame_vm_group_bin_2805 = frame (4k)
frame_vm_group_bin_2806 = frame (4k)
frame_vm_group_bin_2807 = frame (4k)
frame_vm_group_bin_2808 = frame (4k)
frame_vm_group_bin_2809 = frame (4k)
frame_vm_group_bin_2810 = frame (4k)
frame_vm_group_bin_2811 = frame (4k)
frame_vm_group_bin_2812 = frame (4k)
frame_vm_group_bin_2813 = frame (4k)
frame_vm_group_bin_2814 = frame (4k)
frame_vm_group_bin_2815 = frame (4k)
frame_vm_group_bin_2816 = frame (4k)
frame_vm_group_bin_2817 = frame (4k)
frame_vm_group_bin_2818 = frame (4k)
frame_vm_group_bin_2819 = frame (4k)
frame_vm_group_bin_2820 = frame (4k)
frame_vm_group_bin_2821 = frame (4k)
frame_vm_group_bin_2822 = frame (4k)
frame_vm_group_bin_2823 = frame (4k)
frame_vm_group_bin_2824 = frame (4k)
frame_vm_group_bin_2825 = frame (4k)
frame_vm_group_bin_2826 = frame (4k)
frame_vm_group_bin_2827 = frame (4k)
frame_vm_group_bin_2828 = frame (4k)
frame_vm_group_bin_2829 = frame (4k)
frame_vm_group_bin_2830 = frame (4k)
frame_vm_group_bin_2831 = frame (4k)
frame_vm_group_bin_2832 = frame (4k)
frame_vm_group_bin_2833 = frame (4k)
frame_vm_group_bin_2834 = frame (4k)
frame_vm_group_bin_2835 = frame (4k)
frame_vm_group_bin_2836 = frame (4k)
frame_vm_group_bin_2837 = frame (4k)
frame_vm_group_bin_2838 = frame (4k)
frame_vm_group_bin_2839 = frame (4k)
frame_vm_group_bin_2840 = frame (4k)
frame_vm_group_bin_2841 = frame (4k)
frame_vm_group_bin_2842 = frame (4k)
frame_vm_group_bin_2843 = frame (4k)
frame_vm_group_bin_2844 = frame (4k)
frame_vm_group_bin_2845 = frame (4k)
frame_vm_group_bin_2846 = frame (4k)
frame_vm_group_bin_2847 = frame (4k)
frame_vm_group_bin_2848 = frame (4k)
frame_vm_group_bin_2849 = frame (4k)
frame_vm_group_bin_2850 = frame (4k)
frame_vm_group_bin_2851 = frame (4k)
frame_vm_group_bin_2852 = frame (4k)
frame_vm_group_bin_2853 = frame (4k)
frame_vm_group_bin_2854 = frame (4k)
frame_vm_group_bin_2855 = frame (4k)
frame_vm_group_bin_2856 = frame (4k)
frame_vm_group_bin_2857 = frame (4k)
frame_vm_group_bin_2858 = frame (4k)
frame_vm_group_bin_2859 = frame (4k)
frame_vm_group_bin_2860 = frame (4k)
frame_vm_group_bin_2861 = frame (4k)
frame_vm_group_bin_2862 = frame (4k)
frame_vm_group_bin_2863 = frame (4k)
frame_vm_group_bin_2864 = frame (4k)
frame_vm_group_bin_2865 = frame (4k)
frame_vm_group_bin_2866 = frame (4k)
frame_vm_group_bin_2867 = frame (4k)
frame_vm_group_bin_2868 = frame (4k)
frame_vm_group_bin_2869 = frame (4k)
frame_vm_group_bin_2870 = frame (4k)
frame_vm_group_bin_2871 = frame (4k)
frame_vm_group_bin_2872 = frame (4k)
frame_vm_group_bin_2873 = frame (4k)
frame_vm_group_bin_2874 = frame (4k)
frame_vm_group_bin_2875 = frame (4k)
frame_vm_group_bin_2876 = frame (4k)
frame_vm_group_bin_2877 = frame (4k)
frame_vm_group_bin_2878 = frame (4k)
frame_vm_group_bin_2879 = frame (4k)
frame_vm_group_bin_2880 = frame (4k)
frame_vm_group_bin_2881 = frame (4k)
frame_vm_group_bin_2882 = frame (4k)
frame_vm_group_bin_2883 = frame (4k)
frame_vm_group_bin_2884 = frame (4k)
frame_vm_group_bin_2885 = frame (4k)
frame_vm_group_bin_2886 = frame (4k)
frame_vm_group_bin_2887 = frame (4k)
frame_vm_group_bin_2888 = frame (4k)
frame_vm_group_bin_2889 = frame (4k)
frame_vm_group_bin_2890 = frame (4k)
frame_vm_group_bin_2891 = frame (4k)
frame_vm_group_bin_2892 = frame (4k)
frame_vm_group_bin_2893 = frame (4k)
frame_vm_group_bin_2894 = frame (4k)
frame_vm_group_bin_2895 = frame (4k)
frame_vm_group_bin_2896 = frame (4k)
frame_vm_group_bin_2897 = frame (4k)
frame_vm_group_bin_2898 = frame (4k)
frame_vm_group_bin_2899 = frame (4k)
frame_vm_group_bin_2900 = frame (4k)
frame_vm_group_bin_2901 = frame (4k)
frame_vm_group_bin_2902 = frame (4k)
frame_vm_group_bin_2903 = frame (4k)
frame_vm_group_bin_2904 = frame (4k)
frame_vm_group_bin_2905 = frame (4k)
frame_vm_group_bin_2906 = frame (4k)
frame_vm_group_bin_2907 = frame (4k)
frame_vm_group_bin_2908 = frame (4k)
frame_vm_group_bin_2909 = frame (4k)
frame_vm_group_bin_2910 = frame (4k)
frame_vm_group_bin_2911 = frame (4k)
frame_vm_group_bin_2912 = frame (4k)
frame_vm_group_bin_2913 = frame (4k)
frame_vm_group_bin_2914 = frame (4k)
frame_vm_group_bin_2915 = frame (4k)
frame_vm_group_bin_2916 = frame (4k)
frame_vm_group_bin_2917 = frame (4k)
frame_vm_group_bin_2918 = frame (4k)
frame_vm_group_bin_2919 = frame (4k)
frame_vm_group_bin_2920 = frame (4k)
frame_vm_group_bin_2921 = frame (4k)
frame_vm_group_bin_2922 = frame (4k)
frame_vm_group_bin_2923 = frame (4k)
frame_vm_group_bin_2924 = frame (4k)
frame_vm_group_bin_2925 = frame (4k)
frame_vm_group_bin_2926 = frame (4k)
frame_vm_group_bin_2927 = frame (4k)
frame_vm_group_bin_2928 = frame (4k)
frame_vm_group_bin_2929 = frame (4k)
frame_vm_group_bin_2930 = frame (4k)
frame_vm_group_bin_2931 = frame (4k)
frame_vm_group_bin_2932 = frame (4k)
frame_vm_group_bin_2933 = frame (4k)
frame_vm_group_bin_2934 = frame (4k)
frame_vm_group_bin_2935 = frame (4k)
frame_vm_group_bin_2936 = frame (4k)
frame_vm_group_bin_2937 = frame (4k)
frame_vm_group_bin_2938 = frame (4k)
frame_vm_group_bin_2939 = frame (4k)
frame_vm_group_bin_2940 = frame (4k)
frame_vm_group_bin_2941 = frame (4k)
frame_vm_group_bin_2942 = frame (4k)
frame_vm_group_bin_2943 = frame (4k)
frame_vm_group_bin_2944 = frame (4k)
frame_vm_group_bin_2945 = frame (4k)
frame_vm_group_bin_2946 = frame (4k)
frame_vm_group_bin_2947 = frame (4k)
frame_vm_group_bin_2948 = frame (4k)
frame_vm_group_bin_2949 = frame (4k)
frame_vm_group_bin_2950 = frame (4k)
frame_vm_group_bin_2951 = frame (4k)
frame_vm_group_bin_2952 = frame (4k)
frame_vm_group_bin_2953 = frame (4k)
frame_vm_group_bin_2954 = frame (4k)
frame_vm_group_bin_2955 = frame (4k)
frame_vm_group_bin_2956 = frame (4k)
frame_vm_group_bin_2957 = frame (4k)
frame_vm_group_bin_2958 = frame (4k)
frame_vm_group_bin_2959 = frame (4k)
frame_vm_group_bin_2960 = frame (4k)
frame_vm_group_bin_2961 = frame (4k)
frame_vm_group_bin_2962 = frame (4k)
frame_vm_group_bin_2963 = frame (4k)
frame_vm_group_bin_2964 = frame (4k)
frame_vm_group_bin_2965 = frame (4k)
frame_vm_group_bin_2966 = frame (4k)
frame_vm_group_bin_2967 = frame (4k)
frame_vm_group_bin_2968 = frame (4k)
frame_vm_group_bin_2969 = frame (4k)
frame_vm_group_bin_2970 = frame (4k)
frame_vm_group_bin_2971 = frame (4k)
frame_vm_group_bin_2972 = frame (4k)
frame_vm_group_bin_2973 = frame (4k)
frame_vm_group_bin_2974 = frame (4k)
frame_vm_group_bin_2975 = frame (4k)
frame_vm_group_bin_2976 = frame (4k)
frame_vm_group_bin_2977 = frame (4k)
frame_vm_group_bin_2978 = frame (4k)
frame_vm_group_bin_2979 = frame (4k)
frame_vm_group_bin_2980 = frame (4k)
frame_vm_group_bin_2981 = frame (4k)
frame_vm_group_bin_2982 = frame (4k)
frame_vm_group_bin_2983 = frame (4k)
frame_vm_group_bin_2984 = frame (4k)
frame_vm_group_bin_2985 = frame (4k)
frame_vm_group_bin_2986 = frame (4k)
frame_vm_group_bin_2987 = frame (4k)
frame_vm_group_bin_2988 = frame (4k)
frame_vm_group_bin_2989 = frame (4k)
frame_vm_group_bin_2990 = frame (4k)
frame_vm_group_bin_2991 = frame (4k)
frame_vm_group_bin_2992 = frame (4k)
frame_vm_group_bin_2993 = frame (4k)
frame_vm_group_bin_2994 = frame (4k)
frame_vm_group_bin_2995 = frame (4k)
frame_vm_group_bin_2996 = frame (4k)
frame_vm_group_bin_2997 = frame (4k)
frame_vm_group_bin_2998 = frame (4k)
frame_vm_group_bin_2999 = frame (4k)
frame_vm_group_bin_3000 = frame (4k)
frame_vm_group_bin_3001 = frame (4k)
frame_vm_group_bin_3002 = frame (4k)
frame_vm_group_bin_3003 = frame (4k)
frame_vm_group_bin_3004 = frame (4k)
frame_vm_group_bin_3005 = frame (4k)
frame_vm_group_bin_3006 = frame (4k)
frame_vm_group_bin_3007 = frame (4k)
frame_vm_group_bin_3008 = frame (4k)
frame_vm_group_bin_3009 = frame (4k)
frame_vm_group_bin_3010 = frame (4k)
frame_vm_group_bin_3011 = frame (4k)
frame_vm_group_bin_3012 = frame (4k)
frame_vm_group_bin_3013 = frame (4k)
frame_vm_group_bin_3014 = frame (4k)
frame_vm_group_bin_3015 = frame (4k)
frame_vm_group_bin_3016 = frame (4k)
frame_vm_group_bin_3017 = frame (4k)
frame_vm_group_bin_3018 = frame (4k)
frame_vm_group_bin_3019 = frame (4k)
frame_vm_group_bin_3020 = frame (4k)
frame_vm_group_bin_3021 = frame (4k)
frame_vm_group_bin_3022 = frame (4k)
frame_vm_group_bin_3023 = frame (4k)
frame_vm_group_bin_3024 = frame (4k)
frame_vm_group_bin_3025 = frame (4k)
frame_vm_group_bin_3026 = frame (4k)
frame_vm_group_bin_3027 = frame (4k)
frame_vm_group_bin_3028 = frame (4k)
frame_vm_group_bin_3029 = frame (4k)
frame_vm_group_bin_3030 = frame (4k)
frame_vm_group_bin_3031 = frame (4k)
frame_vm_group_bin_3032 = frame (4k)
frame_vm_group_bin_3033 = frame (4k)
frame_vm_group_bin_3034 = frame (4k)
frame_vm_group_bin_3035 = frame (4k)
frame_vm_group_bin_3036 = frame (4k)
frame_vm_group_bin_3037 = frame (4k)
frame_vm_group_bin_3038 = frame (4k)
frame_vm_group_bin_3039 = frame (4k)
frame_vm_group_bin_3040 = frame (4k)
frame_vm_group_bin_3041 = frame (4k)
frame_vm_group_bin_3042 = frame (4k)
frame_vm_group_bin_3043 = frame (4k)
frame_vm_group_bin_3044 = frame (4k)
frame_vm_group_bin_3045 = frame (4k)
frame_vm_group_bin_3046 = frame (4k)
frame_vm_group_bin_3047 = frame (4k)
frame_vm_group_bin_3048 = frame (4k)
frame_vm_group_bin_3049 = frame (4k)
frame_vm_group_bin_3050 = frame (4k)
frame_vm_group_bin_3051 = frame (4k)
frame_vm_group_bin_3052 = frame (4k)
frame_vm_group_bin_3053 = frame (4k)
frame_vm_group_bin_3054 = frame (4k)
frame_vm_group_bin_3055 = frame (4k)
frame_vm_group_bin_3056 = frame (4k)
frame_vm_group_bin_3057 = frame (4k)
frame_vm_group_bin_3058 = frame (4k)
frame_vm_group_bin_3059 = frame (4k)
frame_vm_group_bin_3060 = frame (4k)
frame_vm_group_bin_3061 = frame (4k)
frame_vm_group_bin_3062 = frame (4k)
frame_vm_group_bin_3063 = frame (4k)
frame_vm_group_bin_3064 = frame (4k)
frame_vm_group_bin_3065 = frame (4k)
frame_vm_group_bin_3066 = frame (4k)
frame_vm_group_bin_3067 = frame (4k)
frame_vm_group_bin_3068 = frame (4k)
frame_vm_group_bin_3069 = frame (4k)
frame_vm_group_bin_3070 = frame (4k)
frame_vm_group_bin_3071 = frame (4k)
frame_vm_group_bin_3072 = frame (4k)
frame_vm_group_bin_3073 = frame (4k)
frame_vm_group_bin_3074 = frame (4k)
frame_vm_group_bin_3075 = frame (4k)
frame_vm_group_bin_3076 = frame (4k)
frame_vm_group_bin_3077 = frame (4k)
frame_vm_group_bin_3078 = frame (4k)
frame_vm_group_bin_3079 = frame (4k)
frame_vm_group_bin_3080 = frame (4k)
frame_vm_group_bin_3081 = frame (4k)
frame_vm_group_bin_3082 = frame (4k)
frame_vm_group_bin_3083 = frame (4k)
frame_vm_group_bin_3084 = frame (4k)
frame_vm_group_bin_3085 = frame (4k)
frame_vm_group_bin_3086 = frame (4k)
frame_vm_group_bin_3087 = frame (4k)
frame_vm_group_bin_3088 = frame (4k)
frame_vm_group_bin_3089 = frame (4k)
frame_vm_group_bin_3090 = frame (4k)
frame_vm_group_bin_3091 = frame (4k)
frame_vm_group_bin_3092 = frame (4k)
frame_vm_group_bin_3093 = frame (4k)
frame_vm_group_bin_3094 = frame (4k)
frame_vm_group_bin_3095 = frame (4k)
frame_vm_group_bin_3096 = frame (4k)
frame_vm_group_bin_3097 = frame (4k)
frame_vm_group_bin_3098 = frame (4k)
frame_vm_group_bin_3099 = frame (4k)
frame_vm_group_bin_3100 = frame (4k)
frame_vm_group_bin_3101 = frame (4k)
frame_vm_group_bin_3102 = frame (4k)
frame_vm_group_bin_3103 = frame (4k)
frame_vm_group_bin_3104 = frame (4k)
frame_vm_group_bin_3105 = frame (4k)
frame_vm_group_bin_3106 = frame (4k)
frame_vm_group_bin_3107 = frame (4k)
frame_vm_group_bin_3108 = frame (4k)
frame_vm_group_bin_3109 = frame (4k)
frame_vm_group_bin_3110 = frame (4k)
frame_vm_group_bin_3111 = frame (4k)
frame_vm_group_bin_3112 = frame (4k)
frame_vm_group_bin_3113 = frame (4k)
frame_vm_group_bin_3114 = frame (4k)
frame_vm_group_bin_3115 = frame (4k)
frame_vm_group_bin_3116 = frame (4k)
frame_vm_group_bin_3117 = frame (4k)
frame_vm_group_bin_3118 = frame (4k)
frame_vm_group_bin_3119 = frame (4k)
frame_vm_group_bin_3120 = frame (4k)
frame_vm_group_bin_3121 = frame (4k)
frame_vm_group_bin_3122 = frame (4k)
frame_vm_group_bin_3123 = frame (4k)
frame_vm_group_bin_3124 = frame (4k)
frame_vm_group_bin_3125 = frame (4k)
frame_vm_group_bin_3126 = frame (4k)
frame_vm_group_bin_3127 = frame (4k)
frame_vm_group_bin_3128 = frame (4k)
frame_vm_group_bin_3129 = frame (4k)
frame_vm_group_bin_3130 = frame (4k)
frame_vm_group_bin_3131 = frame (4k)
frame_vm_group_bin_3132 = frame (4k)
frame_vm_group_bin_3133 = frame (4k)
frame_vm_group_bin_3134 = frame (4k)
frame_vm_group_bin_3135 = frame (4k)
frame_vm_group_bin_3136 = frame (4k)
frame_vm_group_bin_3137 = frame (4k)
frame_vm_group_bin_3138 = frame (4k)
frame_vm_group_bin_3139 = frame (4k)
frame_vm_group_bin_3140 = frame (4k)
frame_vm_group_bin_3141 = frame (4k)
frame_vm_group_bin_3142 = frame (4k)
frame_vm_group_bin_3143 = frame (4k)
frame_vm_group_bin_3144 = frame (4k)
frame_vm_group_bin_3145 = frame (4k)
frame_vm_group_bin_3146 = frame (4k)
frame_vm_group_bin_3147 = frame (4k)
frame_vm_group_bin_3148 = frame (4k)
frame_vm_group_bin_3149 = frame (4k)
frame_vm_group_bin_3150 = frame (4k)
frame_vm_group_bin_3151 = frame (4k)
frame_vm_group_bin_3152 = frame (4k)
frame_vm_group_bin_3153 = frame (4k)
frame_vm_group_bin_3154 = frame (4k)
frame_vm_group_bin_3155 = frame (4k)
frame_vm_group_bin_3156 = frame (4k)
frame_vm_group_bin_3157 = frame (4k)
frame_vm_group_bin_3158 = frame (4k)
frame_vm_group_bin_3159 = frame (4k)
frame_vm_group_bin_3160 = frame (4k)
frame_vm_group_bin_3161 = frame (4k)
frame_vm_group_bin_3162 = frame (4k)
frame_vm_group_bin_3163 = frame (4k)
frame_vm_group_bin_3164 = frame (4k)
frame_vm_group_bin_3165 = frame (4k)
frame_vm_group_bin_3166 = frame (4k)
frame_vm_group_bin_3167 = frame (4k)
frame_vm_group_bin_3168 = frame (4k)
frame_vm_group_bin_3169 = frame (4k)
frame_vm_group_bin_3170 = frame (4k)
frame_vm_group_bin_3171 = frame (4k)
frame_vm_group_bin_3172 = frame (4k)
frame_vm_group_bin_3173 = frame (4k)
frame_vm_group_bin_3174 = frame (4k)
frame_vm_group_bin_3175 = frame (4k)
frame_vm_group_bin_3176 = frame (4k)
frame_vm_group_bin_3177 = frame (4k)
frame_vm_group_bin_3178 = frame (4k)
frame_vm_group_bin_3179 = frame (4k)
frame_vm_group_bin_3180 = frame (4k)
frame_vm_group_bin_3181 = frame (4k)
frame_vm_group_bin_3182 = frame (4k)
frame_vm_group_bin_3183 = frame (4k)
frame_vm_group_bin_3184 = frame (4k)
frame_vm_group_bin_3185 = frame (4k)
frame_vm_group_bin_3186 = frame (4k)
frame_vm_group_bin_3187 = frame (4k)
frame_vm_group_bin_3188 = frame (4k)
frame_vm_group_bin_3189 = frame (4k)
frame_vm_group_bin_3190 = frame (4k)
frame_vm_group_bin_3191 = frame (4k)
frame_vm_group_bin_3192 = frame (4k)
frame_vm_group_bin_3193 = frame (4k)
frame_vm_group_bin_3194 = frame (4k)
frame_vm_group_bin_3195 = frame (4k)
frame_vm_group_bin_3196 = frame (4k)
frame_vm_group_bin_3197 = frame (4k)
frame_vm_group_bin_3198 = frame (4k)
frame_vm_group_bin_3199 = frame (4k)
frame_vm_group_bin_3200 = frame (4k)
frame_vm_group_bin_3201 = frame (4k)
frame_vm_group_bin_3202 = frame (4k)
frame_vm_group_bin_3203 = frame (4k)
frame_vm_group_bin_3204 = frame (4k)
frame_vm_group_bin_3205 = frame (4k)
frame_vm_group_bin_3206 = frame (4k)
frame_vm_group_bin_3207 = frame (4k)
frame_vm_group_bin_3208 = frame (4k)
frame_vm_group_bin_3209 = frame (4k)
frame_vm_group_bin_3210 = frame (4k)
frame_vm_group_bin_3211 = frame (4k)
frame_vm_group_bin_3212 = frame (4k)
frame_vm_group_bin_3213 = frame (4k)
frame_vm_group_bin_3214 = frame (4k)
frame_vm_group_bin_3215 = frame (4k)
frame_vm_group_bin_3216 = frame (4k)
frame_vm_group_bin_3217 = frame (4k)
frame_vm_group_bin_3218 = frame (4k)
frame_vm_group_bin_3219 = frame (4k)
frame_vm_group_bin_3220 = frame (4k)
frame_vm_group_bin_3221 = frame (4k)
frame_vm_group_bin_3222 = frame (4k)
frame_vm_group_bin_3223 = frame (4k)
frame_vm_group_bin_3224 = frame (4k)
frame_vm_group_bin_3225 = frame (4k)
frame_vm_group_bin_3226 = frame (4k)
frame_vm_group_bin_3227 = frame (4k)
frame_vm_group_bin_3228 = frame (4k)
frame_vm_group_bin_3229 = frame (4k)
frame_vm_group_bin_3230 = frame (4k)
frame_vm_group_bin_3231 = frame (4k)
frame_vm_group_bin_3232 = frame (4k)
frame_vm_group_bin_3233 = frame (4k)
frame_vm_group_bin_3234 = frame (4k)
frame_vm_group_bin_3235 = frame (4k)
frame_vm_group_bin_3236 = frame (4k)
frame_vm_group_bin_3237 = frame (4k)
frame_vm_group_bin_3238 = frame (4k)
frame_vm_group_bin_3239 = frame (4k)
frame_vm_group_bin_3240 = frame (4k)
frame_vm_group_bin_3241 = frame (4k)
frame_vm_group_bin_3242 = frame (4k)
frame_vm_group_bin_3243 = frame (4k)
frame_vm_group_bin_3244 = frame (4k)
frame_vm_group_bin_3245 = frame (4k)
frame_vm_group_bin_3246 = frame (4k)
frame_vm_group_bin_3247 = frame (4k)
frame_vm_group_bin_3248 = frame (4k)
frame_vm_group_bin_3249 = frame (4k)
frame_vm_group_bin_3250 = frame (4k)
frame_vm_group_bin_3251 = frame (4k)
frame_vm_group_bin_3252 = frame (4k)
frame_vm_group_bin_3253 = frame (4k)
frame_vm_group_bin_3254 = frame (4k)
frame_vm_group_bin_3255 = frame (4k)
frame_vm_group_bin_3256 = frame (4k)
frame_vm_group_bin_3257 = frame (4k)
frame_vm_group_bin_3258 = frame (4k)
frame_vm_group_bin_3259 = frame (4k)
frame_vm_group_bin_3260 = frame (4k)
frame_vm_group_bin_3261 = frame (4k)
frame_vm_group_bin_3262 = frame (4k)
frame_vm_group_bin_3263 = frame (4k)
frame_vm_group_bin_3264 = frame (4k)
frame_vm_group_bin_3265 = frame (4k)
frame_vm_group_bin_3266 = frame (4k)
frame_vm_group_bin_3267 = frame (4k)
frame_vm_group_bin_3268 = frame (4k)
frame_vm_group_bin_3269 = frame (4k)
frame_vm_group_bin_3270 = frame (4k)
frame_vm_group_bin_3271 = frame (4k)
frame_vm_group_bin_3272 = frame (4k)
frame_vm_group_bin_3273 = frame (4k)
frame_vm_group_bin_3274 = frame (4k)
frame_vm_group_bin_3275 = frame (4k)
frame_vm_group_bin_3276 = frame (4k)
frame_vm_group_bin_3277 = frame (4k)
frame_vm_group_bin_3278 = frame (4k)
frame_vm_group_bin_3279 = frame (4k)
frame_vm_group_bin_3280 = frame (4k)
frame_vm_group_bin_3281 = frame (4k)
frame_vm_group_bin_3282 = frame (4k)
frame_vm_group_bin_3283 = frame (4k)
frame_vm_group_bin_3284 = frame (4k)
frame_vm_group_bin_3285 = frame (4k)
frame_vm_group_bin_3286 = frame (4k)
frame_vm_group_bin_3287 = frame (4k)
frame_vm_group_bin_3288 = frame (4k)
frame_vm_group_bin_3289 = frame (4k)
frame_vm_group_bin_3290 = frame (4k)
frame_vm_group_bin_3291 = frame (4k)
frame_vm_group_bin_3292 = frame (4k)
frame_vm_group_bin_3293 = frame (4k)
frame_vm_group_bin_3294 = frame (4k)
frame_vm_group_bin_3295 = frame (4k)
frame_vm_group_bin_3296 = frame (4k)
frame_vm_group_bin_3297 = frame (4k)
frame_vm_group_bin_3298 = frame (4k)
frame_vm_group_bin_3299 = frame (4k)
frame_vm_group_bin_3300 = frame (4k)
frame_vm_group_bin_3301 = frame (4k)
frame_vm_group_bin_3302 = frame (4k)
frame_vm_group_bin_3303 = frame (4k)
frame_vm_group_bin_3304 = frame (4k)
frame_vm_group_bin_3305 = frame (4k)
frame_vm_group_bin_3306 = frame (4k)
frame_vm_group_bin_3307 = frame (4k)
frame_vm_group_bin_3308 = frame (4k)
frame_vm_group_bin_3309 = frame (4k)
frame_vm_group_bin_3310 = frame (4k)
frame_vm_group_bin_3311 = frame (4k)
frame_vm_group_bin_3312 = frame (4k)
frame_vm_group_bin_3313 = frame (4k)
frame_vm_group_bin_3314 = frame (4k)
frame_vm_group_bin_3315 = frame (4k)
frame_vm_group_bin_3316 = frame (4k)
frame_vm_group_bin_3317 = frame (4k)
frame_vm_group_bin_3318 = frame (4k)
frame_vm_group_bin_3319 = frame (4k)
frame_vm_group_bin_3320 = frame (4k)
frame_vm_group_bin_3321 = frame (4k)
frame_vm_group_bin_3322 = frame (4k)
frame_vm_group_bin_3323 = frame (4k)
frame_vm_group_bin_3324 = frame (4k)
frame_vm_group_bin_3325 = frame (4k)
frame_vm_group_bin_3326 = frame (4k)
frame_vm_group_bin_3327 = frame (4k)
frame_vm_group_bin_3328 = frame (4k)
frame_vm_group_bin_3329 = frame (4k)
frame_vm_group_bin_3330 = frame (4k)
frame_vm_group_bin_3331 = frame (4k)
frame_vm_group_bin_3332 = frame (4k)
frame_vm_group_bin_3333 = frame (4k)
frame_vm_group_bin_3334 = frame (4k)
frame_vm_group_bin_3335 = frame (4k)
frame_vm_group_bin_3336 = frame (4k)
frame_vm_group_bin_3337 = frame (4k)
frame_vm_group_bin_3338 = frame (4k)
frame_vm_group_bin_3339 = frame (4k)
frame_vm_group_bin_3340 = frame (4k)
frame_vm_group_bin_3341 = frame (4k)
frame_vm_group_bin_3342 = frame (4k)
frame_vm_group_bin_3343 = frame (4k)
frame_vm_group_bin_3344 = frame (4k)
frame_vm_group_bin_3345 = frame (4k)
frame_vm_group_bin_3346 = frame (4k)
frame_vm_group_bin_3347 = frame (4k)
frame_vm_group_bin_3348 = frame (4k)
frame_vm_group_bin_3349 = frame (4k)
frame_vm_group_bin_3350 = frame (4k)
frame_vm_group_bin_3351 = frame (4k)
frame_vm_group_bin_3352 = frame (4k)
frame_vm_group_bin_3353 = frame (4k)
frame_vm_group_bin_3354 = frame (4k)
frame_vm_group_bin_3355 = frame (4k)
frame_vm_group_bin_3356 = frame (4k)
frame_vm_group_bin_3357 = frame (4k)
frame_vm_group_bin_3358 = frame (4k)
frame_vm_group_bin_3359 = frame (4k)
frame_vm_group_bin_3360 = frame (4k)
frame_vm_group_bin_3361 = frame (4k)
frame_vm_group_bin_3362 = frame (4k)
frame_vm_group_bin_3363 = frame (4k)
frame_vm_group_bin_3364 = frame (4k)
frame_vm_group_bin_3365 = frame (4k)
frame_vm_group_bin_3366 = frame (4k)
frame_vm_group_bin_3367 = frame (4k)
frame_vm_group_bin_3368 = frame (4k)
frame_vm_group_bin_3369 = frame (4k)
frame_vm_group_bin_3370 = frame (4k)
frame_vm_group_bin_3371 = frame (4k)
frame_vm_group_bin_3372 = frame (4k)
frame_vm_group_bin_3373 = frame (4k)
frame_vm_group_bin_3374 = frame (4k)
frame_vm_group_bin_3375 = frame (4k)
frame_vm_group_bin_3376 = frame (4k)
frame_vm_group_bin_3377 = frame (4k)
frame_vm_group_bin_3378 = frame (4k)
frame_vm_group_bin_3379 = frame (4k)
frame_vm_group_bin_3380 = frame (4k)
frame_vm_group_bin_3381 = frame (4k)
frame_vm_group_bin_3382 = frame (4k)
frame_vm_group_bin_3383 = frame (4k)
frame_vm_group_bin_3384 = frame (4k)
frame_vm_group_bin_3385 = frame (4k)
frame_vm_group_bin_3386 = frame (4k)
frame_vm_group_bin_3387 = frame (4k)
frame_vm_group_bin_3388 = frame (4k)
frame_vm_group_bin_3389 = frame (4k)
frame_vm_group_bin_3390 = frame (4k)
frame_vm_group_bin_3391 = frame (4k)
frame_vm_group_bin_3392 = frame (4k)
frame_vm_group_bin_3393 = frame (4k)
frame_vm_group_bin_3394 = frame (4k)
frame_vm_group_bin_3395 = frame (4k)
frame_vm_group_bin_3396 = frame (4k)
frame_vm_group_bin_3397 = frame (4k)
frame_vm_group_bin_3398 = frame (4k)
frame_vm_group_bin_3399 = frame (4k)
frame_vm_group_bin_3400 = frame (4k)
frame_vm_group_bin_3401 = frame (4k)
frame_vm_group_bin_3402 = frame (4k)
frame_vm_group_bin_3403 = frame (4k)
frame_vm_group_bin_3404 = frame (4k)
frame_vm_group_bin_3405 = frame (4k)
frame_vm_group_bin_3406 = frame (4k)
frame_vm_group_bin_3407 = frame (4k)
frame_vm_group_bin_3408 = frame (4k)
frame_vm_group_bin_3409 = frame (4k)
frame_vm_group_bin_3410 = frame (4k)
frame_vm_group_bin_3411 = frame (4k)
frame_vm_group_bin_3412 = frame (4k)
frame_vm_group_bin_3413 = frame (4k)
frame_vm_group_bin_3414 = frame (4k)
frame_vm_group_bin_3415 = frame (4k)
frame_vm_group_bin_3416 = frame (4k)
frame_vm_group_bin_3417 = frame (4k)
frame_vm_group_bin_3418 = frame (4k)
frame_vm_group_bin_3419 = frame (4k)
frame_vm_group_bin_3420 = frame (4k)
frame_vm_group_bin_3421 = frame (4k)
frame_vm_group_bin_3422 = frame (4k)
frame_vm_group_bin_3423 = frame (4k)
frame_vm_group_bin_3424 = frame (4k)
frame_vm_group_bin_3425 = frame (4k)
frame_vm_group_bin_3426 = frame (4k)
frame_vm_group_bin_3427 = frame (4k)
frame_vm_group_bin_3428 = frame (4k)
frame_vm_group_bin_3429 = frame (4k)
frame_vm_group_bin_3430 = frame (4k)
frame_vm_group_bin_3431 = frame (4k)
frame_vm_group_bin_3432 = frame (4k)
frame_vm_group_bin_3433 = frame (4k)
frame_vm_group_bin_3434 = frame (4k)
frame_vm_group_bin_3435 = frame (4k)
frame_vm_group_bin_3436 = frame (4k)
frame_vm_group_bin_3437 = frame (4k)
frame_vm_group_bin_3438 = frame (4k)
frame_vm_group_bin_3439 = frame (4k)
frame_vm_group_bin_3440 = frame (4k)
frame_vm_group_bin_3441 = frame (4k)
frame_vm_group_bin_3442 = frame (4k)
frame_vm_group_bin_3443 = frame (4k)
frame_vm_group_bin_3444 = frame (4k)
frame_vm_group_bin_3445 = frame (4k)
frame_vm_group_bin_3446 = frame (4k)
frame_vm_group_bin_3447 = frame (4k)
frame_vm_group_bin_3448 = frame (4k)
frame_vm_group_bin_3449 = frame (4k)
frame_vm_group_bin_3450 = frame (4k)
frame_vm_group_bin_3451 = frame (4k)
frame_vm_group_bin_3452 = frame (4k)
frame_vm_group_bin_3453 = frame (4k)
frame_vm_group_bin_3454 = frame (4k)
frame_vm_group_bin_3455 = frame (4k)
frame_vm_group_bin_3456 = frame (4k)
frame_vm_group_bin_3457 = frame (4k)
frame_vm_group_bin_3458 = frame (4k)
frame_vm_group_bin_3459 = frame (4k)
frame_vm_group_bin_3460 = frame (4k)
frame_vm_group_bin_3461 = frame (4k)
frame_vm_group_bin_3462 = frame (4k)
frame_vm_group_bin_3463 = frame (4k)
frame_vm_group_bin_3464 = frame (4k)
frame_vm_group_bin_3465 = frame (4k)
frame_vm_group_bin_3466 = frame (4k)
frame_vm_group_bin_3467 = frame (4k)
frame_vm_group_bin_3468 = frame (4k)
frame_vm_group_bin_3469 = frame (4k)
frame_vm_group_bin_3470 = frame (4k)
frame_vm_group_bin_3471 = frame (4k)
frame_vm_group_bin_3472 = frame (4k)
frame_vm_group_bin_3473 = frame (4k)
frame_vm_group_bin_3474 = frame (4k)
frame_vm_group_bin_3475 = frame (4k)
frame_vm_group_bin_3476 = frame (4k)
frame_vm_group_bin_3477 = frame (4k)
frame_vm_group_bin_3478 = frame (4k)
frame_vm_group_bin_3479 = frame (4k)
frame_vm_group_bin_3480 = frame (4k)
frame_vm_group_bin_3481 = frame (4k)
frame_vm_group_bin_3482 = frame (4k)
frame_vm_group_bin_3483 = frame (4k)
frame_vm_group_bin_3484 = frame (4k)
frame_vm_group_bin_3485 = frame (4k)
frame_vm_group_bin_3486 = frame (4k)
frame_vm_group_bin_3487 = frame (4k)
frame_vm_group_bin_3488 = frame (4k)
frame_vm_group_bin_3489 = frame (4k)
frame_vm_group_bin_3490 = frame (4k)
frame_vm_group_bin_3491 = frame (4k)
frame_vm_group_bin_3492 = frame (4k)
frame_vm_group_bin_3493 = frame (4k)
frame_vm_group_bin_3494 = frame (4k)
frame_vm_group_bin_3495 = frame (4k)
frame_vm_group_bin_3496 = frame (4k)
frame_vm_group_bin_3497 = frame (4k)
frame_vm_group_bin_3498 = frame (4k)
frame_vm_group_bin_3499 = frame (4k)
frame_vm_group_bin_3500 = frame (4k)
frame_vm_group_bin_3501 = frame (4k)
frame_vm_group_bin_3502 = frame (4k)
frame_vm_group_bin_3503 = frame (4k)
frame_vm_group_bin_3504 = frame (4k)
frame_vm_group_bin_3505 = frame (4k)
frame_vm_group_bin_3506 = frame (4k)
frame_vm_group_bin_3507 = frame (4k)
frame_vm_group_bin_3508 = frame (4k)
frame_vm_group_bin_3509 = frame (4k)
frame_vm_group_bin_3510 = frame (4k)
frame_vm_group_bin_3511 = frame (4k)
frame_vm_group_bin_3512 = frame (4k)
frame_vm_group_bin_3513 = frame (4k)
frame_vm_group_bin_3514 = frame (4k)
frame_vm_group_bin_3515 = frame (4k)
frame_vm_group_bin_3516 = frame (4k)
frame_vm_group_bin_3517 = frame (4k)
frame_vm_group_bin_3518 = frame (4k)
frame_vm_group_bin_3519 = frame (4k)
frame_vm_group_bin_3520 = frame (4k)
frame_vm_group_bin_3521 = frame (4k)
frame_vm_group_bin_3522 = frame (4k)
frame_vm_group_bin_3523 = frame (4k)
frame_vm_group_bin_3524 = frame (4k)
frame_vm_group_bin_3525 = frame (4k)
frame_vm_group_bin_3526 = frame (4k)
frame_vm_group_bin_3527 = frame (4k)
frame_vm_group_bin_3528 = frame (4k)
frame_vm_group_bin_3529 = frame (4k)
frame_vm_group_bin_3530 = frame (4k)
frame_vm_group_bin_3531 = frame (4k)
frame_vm_group_bin_3532 = frame (4k)
frame_vm_group_bin_3533 = frame (4k)
frame_vm_group_bin_3534 = frame (4k)
frame_vm_group_bin_3535 = frame (4k)
frame_vm_group_bin_3536 = frame (4k)
frame_vm_group_bin_3537 = frame (4k)
frame_vm_group_bin_3538 = frame (4k)
frame_vm_group_bin_3539 = frame (4k)
frame_vm_group_bin_3540 = frame (4k)
frame_vm_group_bin_3541 = frame (4k)
frame_vm_group_bin_3542 = frame (4k)
frame_vm_group_bin_3543 = frame (4k)
frame_vm_group_bin_3544 = frame (4k)
frame_vm_group_bin_3545 = frame (4k)
frame_vm_group_bin_3546 = frame (4k)
frame_vm_group_bin_3547 = frame (4k)
frame_vm_group_bin_3548 = frame (4k)
frame_vm_group_bin_3549 = frame (4k)
frame_vm_group_bin_3550 = frame (4k)
frame_vm_group_bin_3551 = frame (4k)
frame_vm_group_bin_3552 = frame (4k)
frame_vm_group_bin_3553 = frame (4k)
frame_vm_group_bin_3554 = frame (4k)
frame_vm_group_bin_3555 = frame (4k)
frame_vm_group_bin_3556 = frame (4k)
frame_vm_group_bin_3557 = frame (4k)
frame_vm_group_bin_3558 = frame (4k)
frame_vm_group_bin_3559 = frame (4k)
frame_vm_group_bin_3560 = frame (4k)
frame_vm_group_bin_3561 = frame (4k)
frame_vm_group_bin_3562 = frame (4k)
frame_vm_group_bin_3563 = frame (4k)
frame_vm_group_bin_3564 = frame (4k)
frame_vm_group_bin_3565 = frame (4k)
frame_vm_group_bin_3566 = frame (4k)
frame_vm_group_bin_3567 = frame (4k)
frame_vm_group_bin_3568 = frame (4k)
frame_vm_group_bin_3569 = frame (4k)
frame_vm_group_bin_3570 = frame (4k)
frame_vm_group_bin_3571 = frame (4k)
frame_vm_group_bin_3572 = frame (4k)
frame_vm_group_bin_3573 = frame (4k)
frame_vm_group_bin_3574 = frame (4k)
frame_vm_group_bin_3575 = frame (4k)
frame_vm_group_bin_3576 = frame (4k)
frame_vm_group_bin_3577 = frame (4k)
frame_vm_group_bin_3578 = frame (4k)
frame_vm_group_bin_3579 = frame (4k)
frame_vm_group_bin_3580 = frame (4k)
frame_vm_group_bin_3581 = frame (4k)
frame_vm_group_bin_3582 = frame (4k)
frame_vm_group_bin_3583 = frame (4k)
frame_vm_group_bin_3584 = frame (4k)
frame_vm_group_bin_3585 = frame (4k)
frame_vm_group_bin_3586 = frame (4k)
frame_vm_group_bin_3587 = frame (4k)
frame_vm_group_bin_3588 = frame (4k)
frame_vm_group_bin_3589 = frame (4k)
frame_vm_group_bin_3590 = frame (4k)
frame_vm_group_bin_3591 = frame (4k)
frame_vm_group_bin_3592 = frame (4k)
frame_vm_group_bin_3593 = frame (4k)
frame_vm_group_bin_3594 = frame (4k)
frame_vm_group_bin_3595 = frame (4k)
frame_vm_group_bin_3596 = frame (4k)
frame_vm_group_bin_3597 = frame (4k)
frame_vm_group_bin_3598 = frame (4k)
frame_vm_group_bin_3599 = frame (4k)
frame_vm_group_bin_3600 = frame (4k)
frame_vm_group_bin_3601 = frame (4k)
frame_vm_group_bin_3602 = frame (4k)
frame_vm_group_bin_3603 = frame (4k)
frame_vm_group_bin_3604 = frame (4k)
frame_vm_group_bin_3605 = frame (4k)
frame_vm_group_bin_3606 = frame (4k)
frame_vm_group_bin_3607 = frame (4k)
frame_vm_group_bin_3608 = frame (4k)
frame_vm_group_bin_3609 = frame (4k)
frame_vm_group_bin_3610 = frame (4k)
frame_vm_group_bin_3611 = frame (4k)
frame_vm_group_bin_3612 = frame (4k)
frame_vm_group_bin_3613 = frame (4k)
frame_vm_group_bin_3614 = frame (4k)
frame_vm_group_bin_3615 = frame (4k)
frame_vm_group_bin_3616 = frame (4k)
frame_vm_group_bin_3617 = frame (4k)
frame_vm_group_bin_3618 = frame (4k)
frame_vm_group_bin_3619 = frame (4k)
frame_vm_group_bin_3620 = frame (4k)
frame_vm_group_bin_3621 = frame (4k)
frame_vm_group_bin_3622 = frame (4k)
frame_vm_group_bin_3623 = frame (4k)
frame_vm_group_bin_3624 = frame (4k)
frame_vm_group_bin_3625 = frame (4k)
frame_vm_group_bin_3626 = frame (4k)
frame_vm_group_bin_3627 = frame (4k)
frame_vm_group_bin_3628 = frame (4k)
frame_vm_group_bin_3629 = frame (4k)
frame_vm_group_bin_3630 = frame (4k)
frame_vm_group_bin_3631 = frame (4k)
frame_vm_group_bin_3632 = frame (4k)
frame_vm_group_bin_3633 = frame (4k)
frame_vm_group_bin_3634 = frame (4k)
frame_vm_group_bin_3635 = frame (4k)
frame_vm_group_bin_3636 = frame (4k)
frame_vm_group_bin_3637 = frame (4k)
frame_vm_group_bin_3638 = frame (4k)
frame_vm_group_bin_3639 = frame (4k)
frame_vm_group_bin_3640 = frame (4k)
frame_vm_group_bin_3641 = frame (4k)
frame_vm_group_bin_3642 = frame (4k)
frame_vm_group_bin_3643 = frame (4k)
frame_vm_group_bin_3644 = frame (4k)
frame_vm_group_bin_3645 = frame (4k)
frame_vm_group_bin_3646 = frame (4k)
frame_vm_group_bin_3647 = frame (4k)
frame_vm_group_bin_3648 = frame (4k)
frame_vm_group_bin_3649 = frame (4k)
frame_vm_group_bin_3650 = frame (4k)
frame_vm_group_bin_3651 = frame (4k)
frame_vm_group_bin_3652 = frame (4k)
frame_vm_group_bin_3653 = frame (4k)
frame_vm_group_bin_3654 = frame (4k)
frame_vm_group_bin_3655 = frame (4k)
frame_vm_group_bin_3656 = frame (4k)
frame_vm_group_bin_3657 = frame (4k)
frame_vm_group_bin_3658 = frame (4k)
frame_vm_group_bin_3659 = frame (4k)
frame_vm_group_bin_3660 = frame (4k)
frame_vm_group_bin_3661 = frame (4k)
frame_vm_group_bin_3662 = frame (4k)
frame_vm_group_bin_3663 = frame (4k)
frame_vm_group_bin_3664 = frame (4k)
frame_vm_group_bin_3665 = frame (4k)
frame_vm_group_bin_3666 = frame (4k)
frame_vm_group_bin_3667 = frame (4k)
frame_vm_group_bin_3668 = frame (4k)
frame_vm_group_bin_3669 = frame (4k)
frame_vm_group_bin_3670 = frame (4k)
frame_vm_group_bin_3671 = frame (4k)
frame_vm_group_bin_3672 = frame (4k)
frame_vm_group_bin_3673 = frame (4k)
frame_vm_group_bin_3674 = frame (4k)
frame_vm_group_bin_3675 = frame (4k)
frame_vm_group_bin_3676 = frame (4k)
frame_vm_group_bin_3677 = frame (4k)
frame_vm_group_bin_3678 = frame (4k)
frame_vm_group_bin_3679 = frame (4k)
frame_vm_group_bin_3680 = frame (4k)
frame_vm_group_bin_3681 = frame (4k)
frame_vm_group_bin_3682 = frame (4k)
frame_vm_group_bin_3683 = frame (4k)
frame_vm_group_bin_3684 = frame (4k)
frame_vm_group_bin_3685 = frame (4k)
frame_vm_group_bin_3686 = frame (4k)
frame_vm_group_bin_3687 = frame (4k)
frame_vm_group_bin_3688 = frame (4k)
frame_vm_group_bin_3689 = frame (4k)
frame_vm_group_bin_3690 = frame (4k)
frame_vm_group_bin_3691 = frame (4k)
frame_vm_group_bin_3692 = frame (4k)
frame_vm_group_bin_3693 = frame (4k)
frame_vm_group_bin_3694 = frame (4k)
frame_vm_group_bin_3695 = frame (4k)
frame_vm_group_bin_3696 = frame (4k)
frame_vm_group_bin_3697 = frame (4k)
frame_vm_group_bin_3698 = frame (4k)
frame_vm_group_bin_3699 = frame (4k)
frame_vm_group_bin_3700 = frame (4k)
frame_vm_group_bin_3701 = frame (4k)
frame_vm_group_bin_3702 = frame (4k)
frame_vm_group_bin_3703 = frame (4k)
frame_vm_group_bin_3704 = frame (4k)
frame_vm_group_bin_3705 = frame (4k)
frame_vm_group_bin_3706 = frame (4k)
frame_vm_group_bin_3707 = frame (4k)
frame_vm_group_bin_3708 = frame (4k)
frame_vm_group_bin_3709 = frame (4k)
frame_vm_group_bin_3710 = frame (4k)
frame_vm_group_bin_3711 = frame (4k)
frame_vm_group_bin_3712 = frame (4k)
frame_vm_group_bin_3713 = frame (4k)
frame_vm_group_bin_3714 = frame (4k)
frame_vm_group_bin_3715 = frame (4k)
frame_vm_group_bin_3716 = frame (4k)
frame_vm_group_bin_3717 = frame (4k)
frame_vm_group_bin_3718 = frame (4k)
frame_vm_group_bin_3719 = frame (4k)
frame_vm_group_bin_3720 = frame (4k)
frame_vm_group_bin_3721 = frame (4k)
frame_vm_group_bin_3722 = frame (4k)
frame_vm_group_bin_3723 = frame (4k)
frame_vm_group_bin_3724 = frame (4k)
frame_vm_group_bin_3725 = frame (4k)
frame_vm_group_bin_3726 = frame (4k)
frame_vm_group_bin_3727 = frame (4k)
frame_vm_group_bin_3728 = frame (4k)
frame_vm_group_bin_3729 = frame (4k)
frame_vm_group_bin_3730 = frame (4k)
frame_vm_group_bin_3731 = frame (4k)
frame_vm_group_bin_3732 = frame (4k)
frame_vm_group_bin_3733 = frame (4k)
frame_vm_group_bin_3734 = frame (4k)
frame_vm_group_bin_3735 = frame (4k)
frame_vm_group_bin_3736 = frame (4k)
frame_vm_group_bin_3737 = frame (4k)
frame_vm_group_bin_3738 = frame (4k)
frame_vm_group_bin_3739 = frame (4k)
frame_vm_group_bin_3740 = frame (4k)
frame_vm_group_bin_3741 = frame (4k)
frame_vm_group_bin_3742 = frame (4k)
frame_vm_group_bin_3743 = frame (4k)
frame_vm_group_bin_3744 = frame (4k)
frame_vm_group_bin_3745 = frame (4k)
frame_vm_group_bin_3746 = frame (4k)
frame_vm_group_bin_3747 = frame (4k)
frame_vm_group_bin_3748 = frame (4k)
frame_vm_group_bin_3749 = frame (4k)
frame_vm_group_bin_3750 = frame (4k)
frame_vm_group_bin_3751 = frame (4k)
frame_vm_group_bin_3752 = frame (4k)
frame_vm_group_bin_3753 = frame (4k)
frame_vm_group_bin_3754 = frame (4k)
frame_vm_group_bin_3755 = frame (4k)
frame_vm_group_bin_3756 = frame (4k)
frame_vm_group_bin_3757 = frame (4k)
frame_vm_group_bin_3758 = frame (4k)
frame_vm_group_bin_3759 = frame (4k)
frame_vm_group_bin_3760 = frame (4k)
frame_vm_group_bin_3761 = frame (4k)
frame_vm_group_bin_3762 = frame (4k)
frame_vm_group_bin_3763 = frame (4k)
frame_vm_group_bin_3764 = frame (4k)
frame_vm_group_bin_3765 = frame (4k)
frame_vm_group_bin_3766 = frame (4k)
frame_vm_group_bin_3767 = frame (4k)
frame_vm_group_bin_3768 = frame (4k)
frame_vm_group_bin_3769 = frame (4k)
frame_vm_group_bin_3770 = frame (4k)
frame_vm_group_bin_3771 = frame (4k)
frame_vm_group_bin_3772 = frame (4k)
frame_vm_group_bin_3773 = frame (4k)
frame_vm_group_bin_3774 = frame (4k)
frame_vm_group_bin_3775 = frame (4k)
frame_vm_group_bin_3776 = frame (4k)
frame_vm_group_bin_3777 = frame (4k)
frame_vm_group_bin_3778 = frame (4k)
frame_vm_group_bin_3779 = frame (4k)
frame_vm_group_bin_3780 = frame (4k)
frame_vm_group_bin_3781 = frame (4k)
frame_vm_group_bin_3782 = frame (4k)
frame_vm_group_bin_3783 = frame (4k)
frame_vm_group_bin_3784 = frame (4k)
frame_vm_group_bin_3785 = frame (4k)
frame_vm_group_bin_3786 = frame (4k)
frame_vm_group_bin_3787 = frame (4k)
frame_vm_group_bin_3788 = frame (4k)
frame_vm_group_bin_3789 = frame (4k)
frame_vm_group_bin_3790 = frame (4k)
frame_vm_group_bin_3791 = frame (4k)
frame_vm_group_bin_3792 = frame (4k)
frame_vm_group_bin_3793 = frame (4k)
frame_vm_group_bin_3794 = frame (4k)
frame_vm_group_bin_3795 = frame (4k)
frame_vm_group_bin_3796 = frame (4k)
frame_vm_group_bin_3797 = frame (4k)
frame_vm_group_bin_3798 = frame (4k)
frame_vm_group_bin_3799 = frame (4k)
frame_vm_group_bin_3800 = frame (4k)
frame_vm_group_bin_3801 = frame (4k)
frame_vm_group_bin_3802 = frame (4k)
frame_vm_group_bin_3803 = frame (4k)
frame_vm_group_bin_3804 = frame (4k)
frame_vm_group_bin_3805 = frame (4k)
frame_vm_group_bin_3806 = frame (4k)
frame_vm_group_bin_3807 = frame (4k)
frame_vm_group_bin_3808 = frame (4k)
frame_vm_group_bin_3809 = frame (4k)
frame_vm_group_bin_3810 = frame (4k)
frame_vm_group_bin_3811 = frame (4k)
frame_vm_group_bin_3812 = frame (4k)
frame_vm_group_bin_3813 = frame (4k)
frame_vm_group_bin_3814 = frame (4k)
frame_vm_group_bin_3815 = frame (4k)
frame_vm_group_bin_3816 = frame (4k)
frame_vm_group_bin_3817 = frame (4k)
frame_vm_group_bin_3818 = frame (4k)
frame_vm_group_bin_3819 = frame (4k)
frame_vm_group_bin_3820 = frame (4k)
frame_vm_group_bin_3821 = frame (4k)
frame_vm_group_bin_3822 = frame (4k)
frame_vm_group_bin_3823 = frame (4k)
frame_vm_group_bin_3824 = frame (4k)
frame_vm_group_bin_3825 = frame (4k)
frame_vm_group_bin_3826 = frame (4k)
frame_vm_group_bin_3827 = frame (4k)
frame_vm_group_bin_3828 = frame (4k)
frame_vm_group_bin_3829 = frame (4k)
frame_vm_group_bin_3830 = frame (4k)
frame_vm_group_bin_3831 = frame (4k)
frame_vm_group_bin_3832 = frame (4k)
frame_vm_group_bin_3833 = frame (4k)
frame_vm_group_bin_3834 = frame (4k)
frame_vm_group_bin_3835 = frame (4k)
frame_vm_group_bin_3836 = frame (4k)
frame_vm_group_bin_3837 = frame (4k)
frame_vm_group_bin_3838 = frame (4k)
frame_vm_group_bin_3839 = frame (4k)
frame_vm_group_bin_3840 = frame (4k)
frame_vm_group_bin_3841 = frame (4k)
frame_vm_group_bin_3842 = frame (4k)
frame_vm_group_bin_3843 = frame (4k)
frame_vm_group_bin_3844 = frame (4k)
frame_vm_group_bin_3845 = frame (4k)
frame_vm_group_bin_3846 = frame (4k)
frame_vm_group_bin_3847 = frame (4k)
frame_vm_group_bin_3848 = frame (4k)
frame_vm_group_bin_3849 = frame (4k)
frame_vm_group_bin_3850 = frame (4k)
frame_vm_group_bin_3851 = frame (4k)
frame_vm_group_bin_3852 = frame (4k)
frame_vm_group_bin_3853 = frame (4k)
frame_vm_group_bin_3854 = frame (4k)
frame_vm_group_bin_3855 = frame (4k)
frame_vm_group_bin_3856 = frame (4k)
frame_vm_group_bin_3857 = frame (4k)
frame_vm_group_bin_3858 = frame (4k)
frame_vm_group_bin_3859 = frame (4k)
frame_vm_group_bin_3860 = frame (4k)
frame_vm_group_bin_3861 = frame (4k)
frame_vm_group_bin_3862 = frame (4k)
frame_vm_group_bin_3863 = frame (4k)
frame_vm_group_bin_3864 = frame (4k)
frame_vm_group_bin_3865 = frame (4k)
frame_vm_group_bin_3866 = frame (4k)
frame_vm_group_bin_3867 = frame (4k)
frame_vm_group_bin_3868 = frame (4k)
frame_vm_group_bin_3869 = frame (4k)
frame_vm_group_bin_3870 = frame (4k)
frame_vm_group_bin_3871 = frame (4k)
frame_vm_group_bin_3872 = frame (4k)
frame_vm_group_bin_3873 = frame (4k)
frame_vm_group_bin_3874 = frame (4k)
frame_vm_group_bin_3875 = frame (4k)
frame_vm_group_bin_3876 = frame (4k)
frame_vm_group_bin_3877 = frame (4k)
frame_vm_group_bin_3878 = frame (4k)
frame_vm_group_bin_3879 = frame (4k)
frame_vm_group_bin_3880 = frame (4k)
frame_vm_group_bin_3881 = frame (4k)
frame_vm_group_bin_3882 = frame (4k)
frame_vm_group_bin_3883 = frame (4k)
frame_vm_group_bin_3884 = frame (4k)
frame_vm_group_bin_3885 = frame (4k)
frame_vm_group_bin_3886 = frame (4k)
frame_vm_group_bin_3887 = frame (4k)
frame_vm_group_bin_3888 = frame (4k)
frame_vm_group_bin_3889 = frame (4k)
frame_vm_group_bin_3890 = frame (4k)
frame_vm_group_bin_3891 = frame (4k)
frame_vm_group_bin_3892 = frame (4k)
frame_vm_group_bin_3893 = frame (4k)
frame_vm_group_bin_3894 = frame (4k)
frame_vm_group_bin_3895 = frame (4k)
frame_vm_group_bin_3896 = frame (4k)
frame_vm_group_bin_3897 = frame (4k)
frame_vm_group_bin_3898 = frame (4k)
frame_vm_group_bin_3899 = frame (4k)
frame_vm_group_bin_3900 = frame (4k)
frame_vm_group_bin_3901 = frame (4k)
frame_vm_group_bin_3902 = frame (4k)
frame_vm_group_bin_3903 = frame (4k)
frame_vm_group_bin_3904 = frame (4k)
frame_vm_group_bin_3905 = frame (4k)
frame_vm_group_bin_3906 = frame (4k)
frame_vm_group_bin_3907 = frame (4k)
frame_vm_group_bin_3908 = frame (4k)
frame_vm_group_bin_3909 = frame (4k)
frame_vm_group_bin_3910 = frame (4k)
frame_vm_group_bin_3911 = frame (4k)
frame_vm_group_bin_3912 = frame (4k)
frame_vm_group_bin_3913 = frame (4k)
frame_vm_group_bin_3914 = frame (4k)
frame_vm_group_bin_3915 = frame (4k)
frame_vm_group_bin_3916 = frame (4k)
frame_vm_group_bin_3917 = frame (4k)
frame_vm_group_bin_3918 = frame (4k)
frame_vm_group_bin_3919 = frame (4k)
frame_vm_group_bin_3920 = frame (4k)
frame_vm_group_bin_3921 = frame (4k)
frame_vm_group_bin_3922 = frame (4k)
frame_vm_group_bin_3923 = frame (4k)
frame_vm_group_bin_3924 = frame (4k)
frame_vm_group_bin_3925 = frame (4k)
frame_vm_group_bin_3926 = frame (4k)
frame_vm_group_bin_3927 = frame (4k)
frame_vm_group_bin_3928 = frame (4k)
frame_vm_group_bin_3929 = frame (4k)
frame_vm_group_bin_3930 = frame (4k)
frame_vm_group_bin_3931 = frame (4k)
frame_vm_group_bin_3932 = frame (4k)
frame_vm_group_bin_3933 = frame (4k)
frame_vm_group_bin_3934 = frame (4k)
frame_vm_group_bin_3935 = frame (4k)
frame_vm_group_bin_3936 = frame (4k)
frame_vm_group_bin_3937 = frame (4k)
frame_vm_group_bin_3938 = frame (4k)
frame_vm_group_bin_3939 = frame (4k)
frame_vm_group_bin_3940 = frame (4k)
frame_vm_group_bin_3941 = frame (4k)
frame_vm_group_bin_3942 = frame (4k)
frame_vm_group_bin_3943 = frame (4k)
frame_vm_group_bin_3944 = frame (4k)
frame_vm_group_bin_3945 = frame (4k)
frame_vm_group_bin_3946 = frame (4k)
frame_vm_group_bin_3947 = frame (4k)
frame_vm_group_bin_3948 = frame (4k)
frame_vm_group_bin_3949 = frame (4k)
frame_vm_group_bin_3950 = frame (4k)
frame_vm_group_bin_3951 = frame (4k)
frame_vm_group_bin_3952 = frame (4k)
frame_vm_group_bin_3953 = frame (4k)
frame_vm_group_bin_3954 = frame (4k)
frame_vm_group_bin_3955 = frame (4k)
frame_vm_group_bin_3956 = frame (4k)
frame_vm_group_bin_3957 = frame (4k)
frame_vm_group_bin_3958 = frame (4k)
frame_vm_group_bin_3959 = frame (4k)
frame_vm_group_bin_3960 = frame (4k)
frame_vm_group_bin_3961 = frame (4k)
frame_vm_group_bin_3962 = frame (4k)
frame_vm_group_bin_3963 = frame (4k)
frame_vm_group_bin_3964 = frame (4k)
frame_vm_group_bin_3965 = frame (4k)
frame_vm_group_bin_3966 = frame (4k)
frame_vm_group_bin_3967 = frame (4k)
frame_vm_group_bin_3968 = frame (4k)
frame_vm_group_bin_3969 = frame (4k)
frame_vm_group_bin_3970 = frame (4k)
frame_vm_group_bin_3971 = frame (4k)
frame_vm_group_bin_3972 = frame (4k)
frame_vm_group_bin_3973 = frame (4k)
frame_vm_group_bin_3974 = frame (4k)
frame_vm_group_bin_3975 = frame (4k)
frame_vm_group_bin_3976 = frame (4k)
frame_vm_group_bin_3977 = frame (4k)
frame_vm_group_bin_3978 = frame (4k)
frame_vm_group_bin_3979 = frame (4k)
frame_vm_group_bin_3980 = frame (4k)
frame_vm_group_bin_3981 = frame (4k)
frame_vm_group_bin_3982 = frame (4k)
frame_vm_group_bin_3983 = frame (4k)
frame_vm_group_bin_3984 = frame (4k)
frame_vm_group_bin_3985 = frame (4k)
frame_vm_group_bin_3986 = frame (4k)
frame_vm_group_bin_3987 = frame (4k)
frame_vm_group_bin_3988 = frame (4k)
frame_vm_group_bin_3989 = frame (4k)
frame_vm_group_bin_3990 = frame (4k)
frame_vm_group_bin_3991 = frame (4k)
frame_vm_group_bin_3992 = frame (4k)
frame_vm_group_bin_3993 = frame (4k)
frame_vm_group_bin_3994 = frame (4k)
frame_vm_group_bin_3995 = frame (4k)
frame_vm_group_bin_3996 = frame (4k)
frame_vm_group_bin_3997 = frame (4k)
frame_vm_group_bin_3998 = frame (4k)
frame_vm_group_bin_3999 = frame (4k)
frame_vm_group_bin_4000 = frame (4k)
frame_vm_group_bin_4001 = frame (4k)
frame_vm_group_bin_4002 = frame (4k)
frame_vm_group_bin_4003 = frame (4k)
frame_vm_group_bin_4004 = frame (4k)
frame_vm_group_bin_4005 = frame (4k)
frame_vm_group_bin_4006 = frame (4k)
frame_vm_group_bin_4007 = frame (4k)
frame_vm_group_bin_4008 = frame (4k)
frame_vm_group_bin_4009 = frame (4k)
frame_vm_group_bin_4010 = frame (4k)
frame_vm_group_bin_4011 = frame (4k)
frame_vm_group_bin_4012 = frame (4k)
frame_vm_group_bin_4013 = frame (4k)
frame_vm_group_bin_4014 = frame (4k)
frame_vm_group_bin_4015 = frame (4k)
frame_vm_group_bin_4016 = frame (4k)
frame_vm_group_bin_4017 = frame (4k)
frame_vm_group_bin_4018 = frame (4k)
frame_vm_group_bin_4019 = frame (4k)
frame_vm_group_bin_4020 = frame (4k)
frame_vm_group_bin_4021 = frame (4k)
frame_vm_group_bin_4022 = frame (4k)
frame_vm_group_bin_4023 = frame (4k)
frame_vm_group_bin_4024 = frame (4k)
frame_vm_group_bin_4025 = frame (4k)
frame_vm_group_bin_4026 = frame (4k)
frame_vm_group_bin_4027 = frame (4k)
frame_vm_group_bin_4028 = frame (4k)
frame_vm_group_bin_4029 = frame (4k)
frame_vm_group_bin_4030 = frame (4k)
frame_vm_group_bin_4031 = frame (4k)
frame_vm_group_bin_4032 = frame (4k)
frame_vm_group_bin_4033 = frame (4k)
frame_vm_group_bin_4034 = frame (4k)
frame_vm_group_bin_4035 = frame (4k)
frame_vm_group_bin_4036 = frame (4k)
frame_vm_group_bin_4037 = frame (4k)
frame_vm_group_bin_4038 = frame (4k)
frame_vm_group_bin_4039 = frame (4k)
frame_vm_group_bin_4040 = frame (4k)
frame_vm_group_bin_4041 = frame (4k)
frame_vm_group_bin_4042 = frame (4k)
frame_vm_group_bin_4043 = frame (4k)
frame_vm_group_bin_4044 = frame (4k)
frame_vm_group_bin_4045 = frame (4k)
frame_vm_group_bin_4046 = frame (4k)
frame_vm_group_bin_4047 = frame (4k)
frame_vm_group_bin_4048 = frame (4k)
frame_vm_group_bin_4049 = frame (4k)
frame_vm_group_bin_4050 = frame (4k)
frame_vm_group_bin_4051 = frame (4k)
frame_vm_group_bin_4052 = frame (4k)
frame_vm_group_bin_4053 = frame (4k)
frame_vm_group_bin_4054 = frame (4k)
frame_vm_group_bin_4055 = frame (4k)
frame_vm_group_bin_4056 = frame (4k)
frame_vm_group_bin_4057 = frame (4k)
frame_vm_group_bin_4058 = frame (4k)
frame_vm_group_bin_4059 = frame (4k)
frame_vm_group_bin_4060 = frame (4k)
frame_vm_group_bin_4061 = frame (4k)
frame_vm_group_bin_4062 = frame (4k)
frame_vm_group_bin_4063 = frame (4k)
frame_vm_group_bin_4064 = frame (4k)
frame_vm_group_bin_4065 = frame (4k)
frame_vm_group_bin_4066 = frame (4k)
frame_vm_group_bin_4067 = frame (4k)
frame_vm_group_bin_4068 = frame (4k)
frame_vm_group_bin_4069 = frame (4k)
frame_vm_group_bin_4070 = frame (4k)
frame_vm_group_bin_4071 = frame (4k)
frame_vm_group_bin_4072 = frame (4k)
frame_vm_group_bin_4073 = frame (4k)
frame_vm_group_bin_4074 = frame (4k)
frame_vm_group_bin_4075 = frame (4k)
frame_vm_group_bin_4076 = frame (4k)
frame_vm_group_bin_4077 = frame (4k)
frame_vm_group_bin_4078 = frame (4k)
frame_vm_group_bin_4079 = frame (4k)
frame_vm_group_bin_4080 = frame (4k)
frame_vm_group_bin_4081 = frame (4k)
frame_vm_group_bin_4082 = frame (4k)
frame_vm_group_bin_4083 = frame (4k)
frame_vm_group_bin_4084 = frame (4k)
frame_vm_group_bin_4085 = frame (4k)
frame_vm_group_bin_4086 = frame (4k)
frame_vm_group_bin_4087 = frame (4k)
frame_vm_group_bin_4088 = frame (4k)
frame_vm_group_bin_4089 = frame (4k)
frame_vm_group_bin_4090 = frame (4k)
frame_vm_group_bin_4091 = frame (4k)
frame_vm_group_bin_4092 = frame (4k)
frame_vm_group_bin_4093 = frame (4k)
frame_vm_group_bin_4094 = frame (4k)
frame_vm_group_bin_4095 = frame (4k)
frame_vm_group_bin_4096 = frame (4k)
frame_vm_group_bin_4097 = frame (4k)
frame_vm_group_bin_4098 = frame (4k)
frame_vm_group_bin_4099 = frame (4k)
frame_vm_group_bin_4100 = frame (4k)
frame_vm_group_bin_4101 = frame (4k)
frame_vm_group_bin_4102 = frame (4k)
frame_vm_group_bin_4103 = frame (4k)
frame_vm_group_bin_4104 = frame (4k)
frame_vm_group_bin_4105 = frame (4k)
frame_vm_group_bin_4106 = frame (4k)
frame_vm_group_bin_4107 = frame (4k)
frame_vm_group_bin_4108 = frame (4k)
frame_vm_group_bin_4109 = frame (4k)
frame_vm_group_bin_4110 = frame (4k)
frame_vm_group_bin_4111 = frame (4k)
frame_vm_group_bin_4112 = frame (4k)
frame_vm_group_bin_4113 = frame (4k)
frame_vm_group_bin_4114 = frame (4k)
frame_vm_group_bin_4115 = frame (4k)
frame_vm_group_bin_4116 = frame (4k)
frame_vm_group_bin_4117 = frame (4k)
frame_vm_group_bin_4118 = frame (4k)
frame_vm_group_bin_4119 = frame (4k)
frame_vm_group_bin_4120 = frame (4k)
frame_vm_group_bin_4121 = frame (4k)
frame_vm_group_bin_4122 = frame (4k)
frame_vm_group_bin_4123 = frame (4k)
frame_vm_group_bin_4124 = frame (4k)
frame_vm_group_bin_4125 = frame (4k)
frame_vm_group_bin_4126 = frame (4k)
frame_vm_group_bin_4127 = frame (4k)
frame_vm_group_bin_4128 = frame (4k)
frame_vm_group_bin_4129 = frame (4k)
frame_vm_group_bin_4130 = frame (4k)
frame_vm_group_bin_4131 = frame (4k)
frame_vm_group_bin_4132 = frame (4k)
frame_vm_group_bin_4133 = frame (4k)
frame_vm_group_bin_4134 = frame (4k)
frame_vm_group_bin_4135 = frame (4k)
frame_vm_group_bin_4136 = frame (4k)
frame_vm_group_bin_4137 = frame (4k)
frame_vm_group_bin_4138 = frame (4k)
frame_vm_group_bin_4139 = frame (4k)
frame_vm_group_bin_4140 = frame (4k)
frame_vm_group_bin_4141 = frame (4k)
frame_vm_group_bin_4142 = frame (4k)
frame_vm_group_bin_4143 = frame (4k)
frame_vm_group_bin_4144 = frame (4k)
frame_vm_group_bin_4145 = frame (4k)
frame_vm_group_bin_4146 = frame (4k)
frame_vm_group_bin_4147 = frame (4k)
frame_vm_group_bin_4148 = frame (4k)
frame_vm_group_bin_4149 = frame (4k)
frame_vm_group_bin_4150 = frame (4k)
frame_vm_group_bin_4151 = frame (4k)
frame_vm_group_bin_4152 = frame (4k)
frame_vm_group_bin_4153 = frame (4k)
frame_vm_group_bin_4154 = frame (4k)
frame_vm_group_bin_4155 = frame (4k)
frame_vm_group_bin_4156 = frame (4k)
frame_vm_group_bin_4157 = frame (4k)
frame_vm_group_bin_4158 = frame (4k)
frame_vm_group_bin_4159 = frame (4k)
frame_vm_group_bin_4160 = frame (4k)
frame_vm_group_bin_4161 = frame (4k)
frame_vm_group_bin_4162 = frame (4k)
frame_vm_group_bin_4163 = frame (4k)
frame_vm_group_bin_4164 = frame (4k)
frame_vm_group_bin_4165 = frame (4k)
frame_vm_group_bin_4166 = frame (4k)
frame_vm_group_bin_4167 = frame (4k)
frame_vm_group_bin_4168 = frame (4k)
frame_vm_group_bin_4169 = frame (4k)
frame_vm_group_bin_4170 = frame (4k)
frame_vm_group_bin_4171 = frame (4k)
frame_vm_group_bin_4172 = frame (4k)
frame_vm_group_bin_4173 = frame (4k)
frame_vm_group_bin_4174 = frame (4k)
frame_vm_group_bin_4175 = frame (4k)
frame_vm_group_bin_4176 = frame (4k)
frame_vm_group_bin_4177 = frame (4k)
frame_vm_group_bin_4178 = frame (4k)
frame_vm_group_bin_4179 = frame (4k)
frame_vm_group_bin_4180 = frame (4k)
frame_vm_group_bin_4181 = frame (4k)
frame_vm_group_bin_4182 = frame (4k)
frame_vm_group_bin_4183 = frame (4k)
frame_vm_group_bin_4184 = frame (4k)
frame_vm_group_bin_4185 = frame (4k)
frame_vm_group_bin_4186 = frame (4k)
frame_vm_group_bin_4187 = frame (4k)
frame_vm_group_bin_4188 = frame (4k)
frame_vm_group_bin_4189 = frame (4k)
frame_vm_group_bin_4190 = frame (4k)
frame_vm_group_bin_4191 = frame (4k)
frame_vm_group_bin_4192 = frame (4k)
frame_vm_group_bin_4193 = frame (4k)
frame_vm_group_bin_4194 = frame (4k)
frame_vm_group_bin_4195 = frame (4k)
frame_vm_group_bin_4196 = frame (4k)
frame_vm_group_bin_4197 = frame (4k)
frame_vm_group_bin_4198 = frame (4k)
frame_vm_group_bin_4199 = frame (4k)
frame_vm_group_bin_4200 = frame (4k)
frame_vm_group_bin_4201 = frame (4k)
frame_vm_group_bin_4202 = frame (4k)
frame_vm_group_bin_4203 = frame (4k)
frame_vm_group_bin_4204 = frame (4k)
frame_vm_group_bin_4205 = frame (4k)
frame_vm_group_bin_4206 = frame (4k)
frame_vm_group_bin_4207 = frame (4k)
frame_vm_group_bin_4208 = frame (4k)
frame_vm_group_bin_4209 = frame (4k)
frame_vm_group_bin_4210 = frame (4k)
frame_vm_group_bin_4211 = frame (4k)
frame_vm_group_bin_4212 = frame (4k)
frame_vm_group_bin_4213 = frame (4k)
frame_vm_group_bin_4214 = frame (4k)
frame_vm_group_bin_4215 = frame (4k)
frame_vm_group_bin_4216 = frame (4k)
frame_vm_group_bin_4217 = frame (4k)
frame_vm_group_bin_4218 = frame (4k)
frame_vm_group_bin_4219 = frame (4k)
frame_vm_group_bin_4220 = frame (4k)
frame_vm_group_bin_4221 = frame (4k)
frame_vm_group_bin_4222 = frame (4k)
frame_vm_group_bin_4223 = frame (4k)
frame_vm_group_bin_4224 = frame (4k)
frame_vm_group_bin_4225 = frame (4k)
frame_vm_group_bin_4226 = frame (4k)
frame_vm_group_bin_4227 = frame (4k)
frame_vm_group_bin_4228 = frame (4k)
frame_vm_group_bin_4229 = frame (4k)
frame_vm_group_bin_4230 = frame (4k)
frame_vm_group_bin_4231 = frame (4k)
frame_vm_group_bin_4232 = frame (4k)
frame_vm_group_bin_4233 = frame (4k)
frame_vm_group_bin_4234 = frame (4k)
frame_vm_group_bin_4235 = frame (4k)
frame_vm_group_bin_4236 = frame (4k)
frame_vm_group_bin_4237 = frame (4k)
frame_vm_group_bin_4238 = frame (4k)
frame_vm_group_bin_4239 = frame (4k)
frame_vm_group_bin_4240 = frame (4k)
frame_vm_group_bin_4241 = frame (4k)
frame_vm_group_bin_4242 = frame (4k)
frame_vm_group_bin_4243 = frame (4k)
frame_vm_group_bin_4244 = frame (4k)
frame_vm_group_bin_4245 = frame (4k)
frame_vm_group_bin_4246 = frame (4k)
frame_vm_group_bin_4247 = frame (4k)
frame_vm_group_bin_4248 = frame (4k)
frame_vm_group_bin_4249 = frame (4k)
frame_vm_group_bin_4250 = frame (4k)
frame_vm_group_bin_4251 = frame (4k)
frame_vm_group_bin_4252 = frame (4k)
frame_vm_group_bin_4253 = frame (4k)
frame_vm_group_bin_4254 = frame (4k)
frame_vm_group_bin_4255 = frame (4k)
frame_vm_group_bin_4256 = frame (4k)
frame_vm_group_bin_4257 = frame (4k)
frame_vm_group_bin_4258 = frame (4k)
frame_vm_group_bin_4259 = frame (4k)
frame_vm_group_bin_4260 = frame (4k)
frame_vm_group_bin_4261 = frame (4k)
frame_vm_group_bin_4262 = frame (4k)
frame_vm_group_bin_4263 = frame (4k)
frame_vm_group_bin_4264 = frame (4k)
frame_vm_group_bin_4265 = frame (4k)
frame_vm_group_bin_4266 = frame (4k)
frame_vm_group_bin_4267 = frame (4k)
frame_vm_group_bin_4268 = frame (4k)
frame_vm_group_bin_4269 = frame (4k)
frame_vm_group_bin_4270 = frame (4k)
frame_vm_group_bin_4271 = frame (4k)
frame_vm_group_bin_4272 = frame (4k)
frame_vm_group_bin_4273 = frame (4k)
frame_vm_group_bin_4274 = frame (4k)
frame_vm_group_bin_4275 = frame (4k)
frame_vm_group_bin_4276 = frame (4k)
frame_vm_group_bin_4277 = frame (4k)
frame_vm_group_bin_4278 = frame (4k)
frame_vm_group_bin_4279 = frame (4k)
frame_vm_group_bin_4280 = frame (4k)
frame_vm_group_bin_4281 = frame (4k)
frame_vm_group_bin_4282 = frame (4k)
frame_vm_group_bin_4283 = frame (4k)
frame_vm_group_bin_4284 = frame (4k)
frame_vm_group_bin_4285 = frame (4k)
frame_vm_group_bin_4286 = frame (4k)
frame_vm_group_bin_4287 = frame (4k)
frame_vm_group_bin_4288 = frame (4k)
frame_vm_group_bin_4289 = frame (4k)
frame_vm_group_bin_4290 = frame (4k)
frame_vm_group_bin_4291 = frame (4k)
frame_vm_group_bin_4292 = frame (4k)
frame_vm_group_bin_4293 = frame (4k)
frame_vm_group_bin_4294 = frame (4k)
frame_vm_group_bin_4295 = frame (4k)
frame_vm_group_bin_4296 = frame (4k)
frame_vm_group_bin_4297 = frame (4k)
frame_vm_group_bin_4298 = frame (4k)
frame_vm_group_bin_4299 = frame (4k)
frame_vm_group_bin_4300 = frame (4k)
frame_vm_group_bin_4301 = frame (4k)
frame_vm_group_bin_4302 = frame (4k)
frame_vm_group_bin_4303 = frame (4k)
frame_vm_group_bin_4304 = frame (4k)
frame_vm_group_bin_4305 = frame (4k)
frame_vm_group_bin_4306 = frame (4k)
frame_vm_group_bin_4307 = frame (4k)
frame_vm_group_bin_4308 = frame (4k)
frame_vm_group_bin_4309 = frame (4k)
frame_vm_group_bin_4310 = frame (4k)
frame_vm_group_bin_4311 = frame (4k)
frame_vm_group_bin_4312 = frame (4k)
frame_vm_group_bin_4313 = frame (4k)
frame_vm_group_bin_4314 = frame (4k)
frame_vm_group_bin_4315 = frame (4k)
frame_vm_group_bin_4316 = frame (4k)
frame_vm_group_bin_4317 = frame (4k)
frame_vm_group_bin_4318 = frame (4k)
frame_vm_group_bin_4319 = frame (4k)
frame_vm_group_bin_4320 = frame (4k)
frame_vm_group_bin_4321 = frame (4k)
frame_vm_group_bin_4322 = frame (4k)
frame_vm_group_bin_4323 = frame (4k)
frame_vm_group_bin_4324 = frame (4k)
frame_vm_group_bin_4325 = frame (4k)
frame_vm_group_bin_4326 = frame (4k)
frame_vm_group_bin_4327 = frame (4k)
frame_vm_group_bin_4328 = frame (4k)
frame_vm_group_bin_4329 = frame (4k)
frame_vm_group_bin_4330 = frame (4k)
frame_vm_group_bin_4331 = frame (4k)
frame_vm_group_bin_4332 = frame (4k)
frame_vm_group_bin_4333 = frame (4k)
frame_vm_group_bin_4334 = frame (4k)
frame_vm_group_bin_4335 = frame (4k)
frame_vm_group_bin_4336 = frame (4k)
frame_vm_group_bin_4337 = frame (4k)
frame_vm_group_bin_4338 = frame (4k)
frame_vm_group_bin_4339 = frame (4k)
frame_vm_group_bin_4340 = frame (4k)
frame_vm_group_bin_4341 = frame (4k)
frame_vm_group_bin_4342 = frame (4k)
frame_vm_group_bin_4343 = frame (4k)
frame_vm_group_bin_4344 = frame (4k)
frame_vm_group_bin_4345 = frame (4k)
frame_vm_group_bin_4346 = frame (4k)
frame_vm_group_bin_4347 = frame (4k)
frame_vm_group_bin_4348 = frame (4k)
frame_vm_group_bin_4349 = frame (4k)
frame_vm_group_bin_4350 = frame (4k)
frame_vm_group_bin_4351 = frame (4k)
frame_vm_group_bin_4352 = frame (4k)
frame_vm_group_bin_4353 = frame (4k)
frame_vm_group_bin_4354 = frame (4k)
frame_vm_group_bin_4355 = frame (4k)
frame_vm_group_bin_4356 = frame (4k)
frame_vm_group_bin_4357 = frame (4k)
frame_vm_group_bin_4358 = frame (4k)
frame_vm_group_bin_4359 = frame (4k)
frame_vm_group_bin_4360 = frame (4k)
frame_vm_group_bin_4361 = frame (4k)
frame_vm_group_bin_4362 = frame (4k)
frame_vm_group_bin_4363 = frame (4k)
frame_vm_group_bin_4364 = frame (4k)
frame_vm_group_bin_4365 = frame (4k)
frame_vm_group_bin_4366 = frame (4k)
frame_vm_group_bin_4367 = frame (4k)
frame_vm_group_bin_4368 = frame (4k)
frame_vm_group_bin_4369 = frame (4k)
frame_vm_group_bin_4370 = frame (4k)
frame_vm_group_bin_4371 = frame (4k)
frame_vm_group_bin_4372 = frame (4k)
frame_vm_group_bin_4373 = frame (4k)
frame_vm_group_bin_4374 = frame (4k)
frame_vm_group_bin_4375 = frame (4k)
frame_vm_group_bin_4376 = frame (4k)
frame_vm_group_bin_4377 = frame (4k)
frame_vm_group_bin_4378 = frame (4k)
frame_vm_group_bin_4379 = frame (4k)
frame_vm_group_bin_4380 = frame (4k)
frame_vm_group_bin_4381 = frame (4k)
frame_vm_group_bin_4382 = frame (4k)
frame_vm_group_bin_4383 = frame (4k)
frame_vm_group_bin_4384 = frame (4k)
frame_vm_group_bin_4385 = frame (4k)
frame_vm_group_bin_4386 = frame (4k)
frame_vm_group_bin_4387 = frame (4k)
frame_vm_group_bin_4388 = frame (4k)
frame_vm_group_bin_4389 = frame (4k)
frame_vm_group_bin_4390 = frame (4k)
frame_vm_group_bin_4391 = frame (4k)
frame_vm_group_bin_4392 = frame (4k)
frame_vm_group_bin_4393 = frame (4k)
frame_vm_group_bin_4394 = frame (4k)
frame_vm_group_bin_4395 = frame (4k)
frame_vm_group_bin_4396 = frame (4k)
frame_vm_group_bin_4397 = frame (4k)
frame_vm_group_bin_4398 = frame (4k)
frame_vm_group_bin_4399 = frame (4k)
frame_vm_group_bin_4400 = frame (4k)
frame_vm_group_bin_4401 = frame (4k)
frame_vm_group_bin_4402 = frame (4k)
frame_vm_group_bin_4403 = frame (4k)
frame_vm_group_bin_4404 = frame (4k)
frame_vm_group_bin_4405 = frame (4k)
frame_vm_group_bin_4406 = frame (4k)
frame_vm_group_bin_4407 = frame (4k)
frame_vm_group_bin_4408 = frame (4k)
frame_vm_group_bin_4409 = frame (4k)
frame_vm_group_bin_4410 = frame (4k)
frame_vm_group_bin_4411 = frame (4k)
frame_vm_group_bin_4412 = frame (4k)
frame_vm_group_bin_4413 = frame (4k)
frame_vm_group_bin_4414 = frame (4k)
frame_vm_group_bin_4415 = frame (4k)
frame_vm_group_bin_4416 = frame (4k)
frame_vm_group_bin_4417 = frame (4k)
frame_vm_group_bin_4418 = frame (4k)
frame_vm_group_bin_4419 = frame (4k)
frame_vm_group_bin_4420 = frame (4k)
frame_vm_group_bin_4421 = frame (4k)
frame_vm_group_bin_4422 = frame (4k)
frame_vm_group_bin_4423 = frame (4k)
frame_vm_group_bin_4424 = frame (4k)
frame_vm_group_bin_4425 = frame (4k)
frame_vm_group_bin_4426 = frame (4k)
frame_vm_group_bin_4427 = frame (4k)
frame_vm_group_bin_4428 = frame (4k)
frame_vm_group_bin_4429 = frame (4k)
frame_vm_group_bin_4430 = frame (4k)
frame_vm_group_bin_4431 = frame (4k)
frame_vm_group_bin_4432 = frame (4k)
frame_vm_group_bin_4433 = frame (4k)
frame_vm_group_bin_4434 = frame (4k)
frame_vm_group_bin_4435 = frame (4k)
frame_vm_group_bin_4436 = frame (4k)
frame_vm_group_bin_4437 = frame (4k)
frame_vm_group_bin_4438 = frame (4k)
frame_vm_group_bin_4439 = frame (4k)
frame_vm_group_bin_4440 = frame (4k)
frame_vm_group_bin_4441 = frame (4k)
frame_vm_group_bin_4442 = frame (4k)
frame_vm_group_bin_4443 = frame (4k)
frame_vm_group_bin_4444 = frame (4k)
frame_vm_group_bin_4445 = frame (4k)
frame_vm_group_bin_4446 = frame (4k)
frame_vm_group_bin_4447 = frame (4k)
frame_vm_group_bin_4448 = frame (4k)
frame_vm_group_bin_4449 = frame (4k)
frame_vm_group_bin_4450 = frame (4k)
frame_vm_group_bin_4451 = frame (4k)
frame_vm_group_bin_4452 = frame (4k)
frame_vm_group_bin_4453 = frame (4k)
frame_vm_group_bin_4454 = frame (4k)
frame_vm_group_bin_4455 = frame (4k)
frame_vm_group_bin_4456 = frame (4k)
frame_vm_group_bin_4457 = frame (4k)
frame_vm_group_bin_4458 = frame (4k)
frame_vm_group_bin_4459 = frame (4k)
frame_vm_group_bin_4460 = frame (4k)
frame_vm_group_bin_4461 = frame (4k)
frame_vm_group_bin_4462 = frame (4k)
frame_vm_group_bin_4463 = frame (4k)
frame_vm_group_bin_4464 = frame (4k)
frame_vm_group_bin_4465 = frame (4k)
frame_vm_group_bin_4466 = frame (4k)
frame_vm_group_bin_4467 = frame (4k)
frame_vm_group_bin_4468 = frame (4k)
frame_vm_group_bin_4469 = frame (4k)
frame_vm_group_bin_4470 = frame (4k)
frame_vm_group_bin_4471 = frame (4k)
frame_vm_group_bin_4472 = frame (4k)
frame_vm_group_bin_4473 = frame (4k)
frame_vm_group_bin_4474 = frame (4k)
frame_vm_group_bin_4475 = frame (4k)
frame_vm_group_bin_4476 = frame (4k)
frame_vm_group_bin_4477 = frame (4k)
frame_vm_group_bin_4478 = frame (4k)
frame_vm_group_bin_4479 = frame (4k)
frame_vm_group_bin_4480 = frame (4k)
frame_vm_group_bin_4481 = frame (4k)
frame_vm_group_bin_4482 = frame (4k)
frame_vm_group_bin_4483 = frame (4k)
frame_vm_group_bin_4484 = frame (4k)
frame_vm_group_bin_4485 = frame (4k)
frame_vm_group_bin_4486 = frame (4k)
frame_vm_group_bin_4487 = frame (4k)
frame_vm_group_bin_4488 = frame (4k)
frame_vm_group_bin_4489 = frame (4k)
frame_vm_group_bin_4490 = frame (4k)
frame_vm_group_bin_4491 = frame (4k)
frame_vm_group_bin_4492 = frame (4k)
frame_vm_group_bin_4493 = frame (4k)
frame_vm_group_bin_4494 = frame (4k)
frame_vm_group_bin_4495 = frame (4k)
frame_vm_group_bin_4496 = frame (4k)
frame_vm_group_bin_4497 = frame (4k)
frame_vm_group_bin_4498 = frame (4k)
frame_vm_group_bin_4499 = frame (4k)
frame_vm_group_bin_4500 = frame (4k)
frame_vm_group_bin_4501 = frame (4k)
frame_vm_group_bin_4502 = frame (4k)
frame_vm_group_bin_4503 = frame (4k)
frame_vm_group_bin_4504 = frame (4k)
frame_vm_group_bin_4505 = frame (4k)
frame_vm_group_bin_4506 = frame (4k)
frame_vm_group_bin_4507 = frame (4k)
frame_vm_group_bin_4508 = frame (4k)
frame_vm_group_bin_4509 = frame (4k)
frame_vm_group_bin_4510 = frame (4k)
frame_vm_group_bin_4511 = frame (4k)
frame_vm_group_bin_4512 = frame (4k)
frame_vm_group_bin_4513 = frame (4k)
frame_vm_group_bin_4514 = frame (4k)
frame_vm_group_bin_4515 = frame (4k)
frame_vm_group_bin_4516 = frame (4k)
frame_vm_group_bin_4517 = frame (4k)
frame_vm_group_bin_4518 = frame (4k)
frame_vm_group_bin_4519 = frame (4k)
frame_vm_group_bin_4520 = frame (4k)
frame_vm_group_bin_4521 = frame (4k)
frame_vm_group_bin_4522 = frame (4k)
frame_vm_group_bin_4523 = frame (4k)
frame_vm_group_bin_4524 = frame (4k)
frame_vm_group_bin_4525 = frame (4k)
frame_vm_group_bin_4526 = frame (4k)
frame_vm_group_bin_4527 = frame (4k)
frame_vm_group_bin_4528 = frame (4k)
frame_vm_group_bin_4529 = frame (4k)
frame_vm_group_bin_4530 = frame (4k)
frame_vm_group_bin_4531 = frame (4k)
frame_vm_group_bin_4532 = frame (4k)
frame_vm_group_bin_4533 = frame (4k)
frame_vm_group_bin_4534 = frame (4k)
frame_vm_group_bin_4535 = frame (4k)
frame_vm_group_bin_4536 = frame (4k)
frame_vm_group_bin_4537 = frame (4k)
frame_vm_group_bin_4538 = frame (4k)
frame_vm_group_bin_4539 = frame (4k)
frame_vm_group_bin_4540 = frame (4k)
frame_vm_group_bin_4541 = frame (4k)
frame_vm_group_bin_4542 = frame (4k)
frame_vm_group_bin_4543 = frame (4k)
frame_vm_group_bin_4544 = frame (4k)
frame_vm_group_bin_4545 = frame (4k)
frame_vm_group_bin_4546 = frame (4k)
frame_vm_group_bin_4547 = frame (4k)
frame_vm_group_bin_4548 = frame (4k)
frame_vm_group_bin_4549 = frame (4k)
frame_vm_group_bin_4550 = frame (4k)
frame_vm_group_bin_4551 = frame (4k)
frame_vm_group_bin_4552 = frame (4k)
frame_vm_group_bin_4553 = frame (4k)
frame_vm_group_bin_4554 = frame (4k)
frame_vm_group_bin_4555 = frame (4k)
frame_vm_group_bin_4556 = frame (4k)
frame_vm_group_bin_4557 = frame (4k)
frame_vm_group_bin_4558 = frame (4k)
frame_vm_group_bin_4559 = frame (4k)
frame_vm_group_bin_4560 = frame (4k)
frame_vm_group_bin_4561 = frame (4k)
frame_vm_group_bin_4562 = frame (4k)
frame_vm_group_bin_4563 = frame (4k)
frame_vm_group_bin_4564 = frame (4k)
frame_vm_group_bin_4565 = frame (4k)
frame_vm_group_bin_4566 = frame (4k)
frame_vm_group_bin_4567 = frame (4k)
frame_vm_group_bin_4568 = frame (4k)
frame_vm_group_bin_4569 = frame (4k)
frame_vm_group_bin_4570 = frame (4k)
frame_vm_group_bin_4571 = frame (4k)
frame_vm_group_bin_4572 = frame (4k)
frame_vm_group_bin_4573 = frame (4k)
frame_vm_group_bin_4574 = frame (4k)
frame_vm_group_bin_4575 = frame (4k)
frame_vm_group_bin_4576 = frame (4k)
frame_vm_group_bin_4577 = frame (4k)
frame_vm_group_bin_4578 = frame (4k)
frame_vm_group_bin_4579 = frame (4k)
frame_vm_group_bin_4580 = frame (4k)
frame_vm_group_bin_4581 = frame (4k)
frame_vm_group_bin_4582 = frame (4k)
frame_vm_group_bin_4583 = frame (4k)
frame_vm_group_bin_4584 = frame (4k)
frame_vm_group_bin_4585 = frame (4k)
frame_vm_group_bin_4586 = frame (4k)
frame_vm_group_bin_4587 = frame (4k)
frame_vm_group_bin_4588 = frame (4k)
frame_vm_group_bin_4589 = frame (4k)
frame_vm_group_bin_4590 = frame (4k)
frame_vm_group_bin_4591 = frame (4k)
frame_vm_group_bin_4592 = frame (4k)
frame_vm_group_bin_4593 = frame (4k)
frame_vm_group_bin_4594 = frame (4k)
frame_vm_group_bin_4595 = frame (4k)
frame_vm_group_bin_4596 = frame (4k)
frame_vm_group_bin_4597 = frame (4k)
frame_vm_group_bin_4598 = frame (4k)
frame_vm_group_bin_4599 = frame (4k)
frame_vm_group_bin_4600 = frame (4k)
frame_vm_group_bin_4601 = frame (4k)
frame_vm_group_bin_4602 = frame (4k)
frame_vm_group_bin_4603 = frame (4k)
frame_vm_group_bin_4604 = frame (4k)
frame_vm_group_bin_4605 = frame (4k)
frame_vm_group_bin_4606 = frame (4k)
frame_vm_group_bin_4607 = frame (4k)
frame_vm_group_bin_4608 = frame (4k)
frame_vm_group_bin_4609 = frame (4k)
frame_vm_group_bin_4610 = frame (4k)
frame_vm_group_bin_4611 = frame (4k)
frame_vm_group_bin_4612 = frame (4k)
frame_vm_group_bin_4613 = frame (4k)
frame_vm_group_bin_4614 = frame (4k)
frame_vm_group_bin_4615 = frame (4k)
frame_vm_group_bin_4616 = frame (4k)
frame_vm_group_bin_4617 = frame (4k)
frame_vm_group_bin_4618 = frame (4k)
frame_vm_group_bin_4619 = frame (4k)
frame_vm_group_bin_4620 = frame (4k)
frame_vm_group_bin_4621 = frame (4k)
frame_vm_group_bin_4622 = frame (4k)
frame_vm_group_bin_4623 = frame (4k)
frame_vm_group_bin_4624 = frame (4k)
frame_vm_group_bin_4625 = frame (4k)
frame_vm_group_bin_4626 = frame (4k)
frame_vm_group_bin_4627 = frame (4k)
frame_vm_group_bin_4628 = frame (4k)
frame_vm_group_bin_4629 = frame (4k)
frame_vm_group_bin_4630 = frame (4k)
frame_vm_group_bin_4631 = frame (4k)
frame_vm_group_bin_4632 = frame (4k)
frame_vm_group_bin_4633 = frame (4k)
frame_vm_group_bin_4634 = frame (4k)
frame_vm_group_bin_4635 = frame (4k)
frame_vm_group_bin_4636 = frame (4k)
frame_vm_group_bin_4637 = frame (4k)
frame_vm_group_bin_4638 = frame (4k)
frame_vm_group_bin_4639 = frame (4k)
frame_vm_group_bin_4640 = frame (4k)
frame_vm_group_bin_4641 = frame (4k)
frame_vm_group_bin_4642 = frame (4k)
frame_vm_group_bin_4643 = frame (4k)
frame_vm_group_bin_4644 = frame (4k)
frame_vm_group_bin_4645 = frame (4k)
frame_vm_group_bin_4646 = frame (4k)
frame_vm_group_bin_4647 = frame (4k)
frame_vm_group_bin_4648 = frame (4k)
frame_vm_group_bin_4649 = frame (4k)
frame_vm_group_bin_4650 = frame (4k)
frame_vm_group_bin_4651 = frame (4k)
frame_vm_group_bin_4652 = frame (4k)
frame_vm_group_bin_4653 = frame (4k)
frame_vm_group_bin_4654 = frame (4k)
frame_vm_group_bin_4655 = frame (4k)
frame_vm_group_bin_4656 = frame (4k)
frame_vm_group_bin_4657 = frame (4k)
frame_vm_group_bin_4658 = frame (4k)
frame_vm_group_bin_4659 = frame (4k)
frame_vm_group_bin_4660 = frame (4k)
frame_vm_group_bin_4661 = frame (4k)
frame_vm_group_bin_4662 = frame (4k)
frame_vm_group_bin_4663 = frame (4k)
frame_vm_group_bin_4664 = frame (4k)
frame_vm_group_bin_4665 = frame (4k)
frame_vm_group_bin_4666 = frame (4k)
frame_vm_group_bin_4667 = frame (4k)
frame_vm_group_bin_4668 = frame (4k)
frame_vm_group_bin_4669 = frame (4k)
frame_vm_group_bin_4670 = frame (4k)
frame_vm_group_bin_4671 = frame (4k)
frame_vm_group_bin_4672 = frame (4k)
frame_vm_group_bin_4673 = frame (4k)
frame_vm_group_bin_4674 = frame (4k)
frame_vm_group_bin_4675 = frame (4k)
frame_vm_group_bin_4676 = frame (4k)
frame_vm_group_bin_4677 = frame (4k)
frame_vm_group_bin_4678 = frame (4k)
frame_vm_group_bin_4679 = frame (4k)
frame_vm_group_bin_4680 = frame (4k)
frame_vm_group_bin_4681 = frame (4k)
frame_vm_group_bin_4682 = frame (4k)
frame_vm_group_bin_4683 = frame (4k)
frame_vm_group_bin_4684 = frame (4k)
frame_vm_group_bin_4685 = frame (4k)
frame_vm_group_bin_4686 = frame (4k)
frame_vm_group_bin_4687 = frame (4k)
frame_vm_group_bin_4688 = frame (4k)
frame_vm_group_bin_4689 = frame (4k)
frame_vm_group_bin_4690 = frame (4k)
frame_vm_group_bin_4691 = frame (4k)
frame_vm_group_bin_4692 = frame (4k)
frame_vm_group_bin_4693 = frame (4k)
frame_vm_group_bin_4694 = frame (4k)
frame_vm_group_bin_4695 = frame (4k)
frame_vm_group_bin_4696 = frame (4k)
frame_vm_group_bin_4697 = frame (4k)
frame_vm_group_bin_4698 = frame (4k)
frame_vm_group_bin_4699 = frame (4k)
frame_vm_group_bin_4700 = frame (4k)
frame_vm_group_bin_4701 = frame (4k)
frame_vm_group_bin_4702 = frame (4k)
frame_vm_group_bin_4703 = frame (4k)
frame_vm_group_bin_4704 = frame (4k)
frame_vm_group_bin_4705 = frame (4k)
frame_vm_group_bin_4706 = frame (4k)
frame_vm_group_bin_4707 = frame (4k)
frame_vm_group_bin_4708 = frame (4k)
frame_vm_group_bin_4709 = frame (4k)
frame_vm_group_bin_4710 = frame (4k)
frame_vm_group_bin_4711 = frame (4k)
frame_vm_group_bin_4712 = frame (4k)
frame_vm_group_bin_4713 = frame (4k)
frame_vm_group_bin_4714 = frame (4k)
frame_vm_group_bin_4715 = frame (4k)
frame_vm_group_bin_4716 = frame (4k)
frame_vm_group_bin_4717 = frame (4k)
frame_vm_group_bin_4718 = frame (4k)
frame_vm_group_bin_4719 = frame (4k)
frame_vm_group_bin_4720 = frame (4k)
frame_vm_group_bin_4721 = frame (4k)
frame_vm_group_bin_4722 = frame (4k)
frame_vm_group_bin_4723 = frame (4k)
frame_vm_group_bin_4724 = frame (4k)
frame_vm_group_bin_4725 = frame (4k)
frame_vm_group_bin_4726 = frame (4k)
frame_vm_group_bin_4727 = frame (4k)
frame_vm_group_bin_4728 = frame (4k)
frame_vm_group_bin_4729 = frame (4k)
frame_vm_group_bin_4730 = frame (4k)
frame_vm_group_bin_4731 = frame (4k)
frame_vm_group_bin_4732 = frame (4k)
frame_vm_group_bin_4733 = frame (4k)
frame_vm_group_bin_4734 = frame (4k)
frame_vm_group_bin_4735 = frame (4k)
frame_vm_group_bin_4736 = frame (4k)
frame_vm_group_bin_4737 = frame (4k)
frame_vm_group_bin_4738 = frame (4k)
frame_vm_group_bin_4739 = frame (4k)
frame_vm_group_bin_4740 = frame (4k)
frame_vm_group_bin_4741 = frame (4k)
frame_vm_group_bin_4742 = frame (4k)
frame_vm_group_bin_4743 = frame (4k)
frame_vm_group_bin_4744 = frame (4k)
frame_vm_group_bin_4745 = frame (4k)
frame_vm_group_bin_4746 = frame (4k)
frame_vm_group_bin_4747 = frame (4k)
frame_vm_group_bin_4748 = frame (4k)
frame_vm_group_bin_4749 = frame (4k)
frame_vm_group_bin_4750 = frame (4k)
frame_vm_group_bin_4751 = frame (4k)
frame_vm_group_bin_4752 = frame (4k)
frame_vm_group_bin_4753 = frame (4k)
frame_vm_group_bin_4754 = frame (4k)
frame_vm_group_bin_4755 = frame (4k)
frame_vm_group_bin_4756 = frame (4k)
frame_vm_group_bin_4757 = frame (4k)
frame_vm_group_bin_4758 = frame (4k)
frame_vm_group_bin_4759 = frame (4k)
frame_vm_group_bin_4760 = frame (4k)
frame_vm_group_bin_4761 = frame (4k)
frame_vm_group_bin_4762 = frame (4k)
frame_vm_group_bin_4763 = frame (4k)
frame_vm_group_bin_4764 = frame (4k)
frame_vm_group_bin_4765 = frame (4k)
frame_vm_group_bin_4766 = frame (4k)
frame_vm_group_bin_4767 = frame (4k)
frame_vm_group_bin_4768 = frame (4k)
frame_vm_group_bin_4769 = frame (4k)
frame_vm_group_bin_4770 = frame (4k)
frame_vm_group_bin_4771 = frame (4k)
frame_vm_group_bin_4772 = frame (4k)
frame_vm_group_bin_4773 = frame (4k)
frame_vm_group_bin_4774 = frame (4k)
frame_vm_group_bin_4775 = frame (4k)
frame_vm_group_bin_4776 = frame (4k)
frame_vm_group_bin_4777 = frame (4k)
frame_vm_group_bin_4778 = frame (4k)
frame_vm_group_bin_4779 = frame (4k)
frame_vm_group_bin_4780 = frame (4k)
frame_vm_group_bin_4781 = frame (4k)
frame_vm_group_bin_4782 = frame (4k)
frame_vm_group_bin_4783 = frame (4k)
frame_vm_group_bin_4784 = frame (4k)
frame_vm_group_bin_4785 = frame (4k)
frame_vm_group_bin_4786 = frame (4k)
frame_vm_group_bin_4787 = frame (4k)
frame_vm_group_bin_4788 = frame (4k)
frame_vm_group_bin_4789 = frame (4k)
frame_vm_group_bin_4790 = frame (4k)
frame_vm_group_bin_4791 = frame (4k)
frame_vm_group_bin_4792 = frame (4k)
frame_vm_group_bin_4793 = frame (4k)
frame_vm_group_bin_4794 = frame (4k)
frame_vm_group_bin_4795 = frame (4k)
frame_vm_group_bin_4796 = frame (4k)
frame_vm_group_bin_4797 = frame (4k)
frame_vm_group_bin_4798 = frame (4k)
frame_vm_group_bin_4799 = frame (4k)
frame_vm_group_bin_4800 = frame (4k)
frame_vm_group_bin_4801 = frame (4k)
frame_vm_group_bin_4802 = frame (4k)
frame_vm_group_bin_4803 = frame (4k)
frame_vm_group_bin_4804 = frame (4k)
frame_vm_group_bin_4805 = frame (4k)
frame_vm_group_bin_4806 = frame (4k)
frame_vm_group_bin_4807 = frame (4k)
frame_vm_group_bin_4808 = frame (4k)
frame_vm_group_bin_4809 = frame (4k)
frame_vm_group_bin_4810 = frame (4k)
frame_vm_group_bin_4811 = frame (4k)
frame_vm_group_bin_4812 = frame (4k)
frame_vm_group_bin_4813 = frame (4k)
frame_vm_group_bin_4814 = frame (4k)
frame_vm_group_bin_4815 = frame (4k)
frame_vm_group_bin_4816 = frame (4k)
frame_vm_group_bin_4817 = frame (4k)
frame_vm_group_bin_4818 = frame (4k)
frame_vm_group_bin_4819 = frame (4k)
frame_vm_group_bin_4820 = frame (4k)
frame_vm_group_bin_4821 = frame (4k)
frame_vm_group_bin_4822 = frame (4k)
frame_vm_group_bin_4823 = frame (4k)
frame_vm_group_bin_4824 = frame (4k)
frame_vm_group_bin_4825 = frame (4k)
frame_vm_group_bin_4826 = frame (4k)
frame_vm_group_bin_4827 = frame (4k)
frame_vm_group_bin_4828 = frame (4k)
frame_vm_group_bin_4829 = frame (4k)
frame_vm_group_bin_4830 = frame (4k)
frame_vm_group_bin_4831 = frame (4k)
frame_vm_group_bin_4832 = frame (4k)
frame_vm_group_bin_4833 = frame (4k)
frame_vm_group_bin_4834 = frame (4k)
frame_vm_group_bin_4835 = frame (4k)
frame_vm_group_bin_4836 = frame (4k)
frame_vm_group_bin_4837 = frame (4k)
frame_vm_group_bin_4838 = frame (4k)
frame_vm_group_bin_4839 = frame (4k)
frame_vm_group_bin_4840 = frame (4k)
frame_vm_group_bin_4841 = frame (4k)
frame_vm_group_bin_4842 = frame (4k)
frame_vm_group_bin_4843 = frame (4k)
frame_vm_group_bin_4844 = frame (4k)
frame_vm_group_bin_4845 = frame (4k)
frame_vm_group_bin_4846 = frame (4k)
frame_vm_group_bin_4847 = frame (4k)
frame_vm_group_bin_4848 = frame (4k)
frame_vm_group_bin_4849 = frame (4k)
frame_vm_group_bin_4850 = frame (4k)
frame_vm_group_bin_4851 = frame (4k)
frame_vm_group_bin_4852 = frame (4k)
frame_vm_group_bin_4853 = frame (4k)
frame_vm_group_bin_4854 = frame (4k)
frame_vm_group_bin_4855 = frame (4k)
frame_vm_group_bin_4856 = frame (4k)
frame_vm_group_bin_4857 = frame (4k)
frame_vm_group_bin_4858 = frame (4k)
frame_vm_group_bin_4859 = frame (4k)
frame_vm_group_bin_4860 = frame (4k)
frame_vm_group_bin_4861 = frame (4k)
frame_vm_group_bin_4862 = frame (4k)
frame_vm_group_bin_4863 = frame (4k)
frame_vm_group_bin_4864 = frame (4k)
frame_vm_group_bin_4865 = frame (4k)
frame_vm_group_bin_4866 = frame (4k)
frame_vm_group_bin_4867 = frame (4k)
frame_vm_group_bin_4868 = frame (4k)
frame_vm_group_bin_4869 = frame (4k)
frame_vm_group_bin_4870 = frame (4k)
frame_vm_group_bin_4871 = frame (4k)
frame_vm_group_bin_4872 = frame (4k)
frame_vm_group_bin_4873 = frame (4k)
frame_vm_group_bin_4874 = frame (4k)
frame_vm_group_bin_4875 = frame (4k)
frame_vm_group_bin_4876 = frame (4k)
frame_vm_group_bin_4877 = frame (4k)
frame_vm_group_bin_4878 = frame (4k)
frame_vm_group_bin_4879 = frame (4k)
frame_vm_group_bin_4880 = frame (4k)
frame_vm_group_bin_4881 = frame (4k)
frame_vm_group_bin_4882 = frame (4k)
frame_vm_group_bin_4883 = frame (4k)
frame_vm_group_bin_4884 = frame (4k)
frame_vm_group_bin_4885 = frame (4k)
frame_vm_group_bin_4886 = frame (4k)
frame_vm_group_bin_4887 = frame (4k)
frame_vm_group_bin_4888 = frame (4k)
frame_vm_group_bin_4889 = frame (4k)
frame_vm_group_bin_4890 = frame (4k)
frame_vm_group_bin_4891 = frame (4k)
frame_vm_group_bin_4892 = frame (4k)
frame_vm_group_bin_4893 = frame (4k)
frame_vm_group_bin_4894 = frame (4k)
frame_vm_group_bin_4895 = frame (4k)
frame_vm_group_bin_4896 = frame (4k)
frame_vm_group_bin_4897 = frame (4k)
frame_vm_group_bin_4898 = frame (4k)
frame_vm_group_bin_4899 = frame (4k)
frame_vm_group_bin_4900 = frame (4k)
frame_vm_group_bin_4901 = frame (4k)
frame_vm_group_bin_4902 = frame (4k)
frame_vm_group_bin_4903 = frame (4k)
frame_vm_group_bin_4904 = frame (4k)
frame_vm_group_bin_4905 = frame (4k)
frame_vm_group_bin_4906 = frame (4k)
frame_vm_group_bin_4907 = frame (4k)
frame_vm_group_bin_4908 = frame (4k)
frame_vm_group_bin_4909 = frame (4k)
frame_vm_group_bin_4910 = frame (4k)
frame_vm_group_bin_4911 = frame (4k)
frame_vm_group_bin_4912 = frame (4k)
frame_vm_group_bin_4913 = frame (4k)
frame_vm_group_bin_4914 = frame (4k)
frame_vm_group_bin_4915 = frame (4k)
frame_vm_group_bin_4916 = frame (4k)
frame_vm_group_bin_4917 = frame (4k)
frame_vm_group_bin_4918 = frame (4k)
frame_vm_group_bin_4919 = frame (4k)
frame_vm_group_bin_4920 = frame (4k)
frame_vm_group_bin_4921 = frame (4k)
frame_vm_group_bin_4922 = frame (4k)
frame_vm_group_bin_4923 = frame (4k)
frame_vm_group_bin_4924 = frame (4k)
frame_vm_group_bin_4925 = frame (4k)
frame_vm_group_bin_4926 = frame (4k)
frame_vm_group_bin_4927 = frame (4k)
frame_vm_group_bin_4928 = frame (4k)
frame_vm_group_bin_4929 = frame (4k)
frame_vm_group_bin_4930 = frame (4k)
frame_vm_group_bin_4931 = frame (4k)
frame_vm_group_bin_4932 = frame (4k)
frame_vm_group_bin_4933 = frame (4k)
frame_vm_group_bin_4934 = frame (4k)
frame_vm_group_bin_4935 = frame (4k)
frame_vm_group_bin_4936 = frame (4k)
frame_vm_group_bin_4937 = frame (4k)
frame_vm_group_bin_4938 = frame (4k)
frame_vm_group_bin_4939 = frame (4k)
frame_vm_group_bin_4940 = frame (4k)
frame_vm_group_bin_4941 = frame (4k)
frame_vm_group_bin_4942 = frame (4k)
frame_vm_group_bin_4943 = frame (4k)
frame_vm_group_bin_4944 = frame (4k)
frame_vm_group_bin_4945 = frame (4k)
frame_vm_group_bin_4946 = frame (4k)
frame_vm_group_bin_4947 = frame (4k)
frame_vm_group_bin_4948 = frame (4k)
frame_vm_group_bin_4949 = frame (4k)
frame_vm_group_bin_4950 = frame (4k)
frame_vm_group_bin_4951 = frame (4k)
frame_vm_group_bin_4952 = frame (4k)
frame_vm_group_bin_4953 = frame (4k)
frame_vm_group_bin_4954 = frame (4k)
frame_vm_group_bin_4955 = frame (4k)
frame_vm_group_bin_4956 = frame (4k)
frame_vm_group_bin_4957 = frame (4k)
frame_vm_group_bin_4958 = frame (4k)
frame_vm_group_bin_4959 = frame (4k)
frame_vm_group_bin_4960 = frame (4k)
frame_vm_group_bin_4961 = frame (4k)
frame_vm_group_bin_4962 = frame (4k)
frame_vm_group_bin_4963 = frame (4k)
frame_vm_group_bin_4964 = frame (4k)
frame_vm_group_bin_4965 = frame (4k)
frame_vm_group_bin_4966 = frame (4k)
frame_vm_group_bin_4967 = frame (4k)
frame_vm_group_bin_4968 = frame (4k)
frame_vm_group_bin_4969 = frame (4k)
frame_vm_group_bin_4970 = frame (4k)
frame_vm_group_bin_4971 = frame (4k)
frame_vm_group_bin_4972 = frame (4k)
frame_vm_group_bin_4973 = frame (4k)
frame_vm_group_bin_4974 = frame (4k)
frame_vm_group_bin_4975 = frame (4k)
frame_vm_group_bin_4976 = frame (4k)
frame_vm_group_bin_4977 = frame (4k)
frame_vm_group_bin_4978 = frame (4k)
frame_vm_group_bin_4979 = frame (4k)
frame_vm_group_bin_4980 = frame (4k)
frame_vm_group_bin_4981 = frame (4k)
frame_vm_group_bin_4982 = frame (4k)
frame_vm_group_bin_4983 = frame (4k)
frame_vm_group_bin_4984 = frame (4k)
frame_vm_group_bin_4985 = frame (4k)
frame_vm_group_bin_4986 = frame (4k)
frame_vm_group_bin_4987 = frame (4k)
frame_vm_group_bin_4988 = frame (4k)
frame_vm_group_bin_4989 = frame (4k)
frame_vm_group_bin_4990 = frame (4k)
frame_vm_group_bin_4991 = frame (4k)
frame_vm_group_bin_4992 = frame (4k)
frame_vm_group_bin_4993 = frame (4k)
frame_vm_group_bin_4994 = frame (4k)
frame_vm_group_bin_4995 = frame (4k)
frame_vm_group_bin_4996 = frame (4k)
frame_vm_group_bin_4997 = frame (4k)
frame_vm_group_bin_4998 = frame (4k)
frame_vm_group_bin_4999 = frame (4k)
frame_vm_group_bin_5000 = frame (4k)
frame_vm_group_bin_5001 = frame (4k)
frame_vm_group_bin_5002 = frame (4k)
frame_vm_group_bin_5003 = frame (4k)
frame_vm_group_bin_5004 = frame (4k)
frame_vm_group_bin_5005 = frame (4k)
frame_vm_group_bin_5006 = frame (4k)
frame_vm_group_bin_5007 = frame (4k)
frame_vm_group_bin_5008 = frame (4k)
frame_vm_group_bin_5009 = frame (4k)
frame_vm_group_bin_5010 = frame (4k)
frame_vm_group_bin_5011 = frame (4k)
frame_vm_group_bin_5012 = frame (4k)
frame_vm_group_bin_5013 = frame (4k)
frame_vm_group_bin_5014 = frame (4k)
frame_vm_group_bin_5015 = frame (4k)
frame_vm_group_bin_5016 = frame (4k)
frame_vm_group_bin_5017 = frame (4k)
frame_vm_group_bin_5018 = frame (4k)
frame_vm_group_bin_5019 = frame (4k)
frame_vm_group_bin_5020 = frame (4k)
frame_vm_group_bin_5021 = frame (4k)
frame_vm_group_bin_5022 = frame (4k)
frame_vm_group_bin_5023 = frame (4k)
frame_vm_group_bin_5024 = frame (4k)
frame_vm_group_bin_5025 = frame (4k)
frame_vm_group_bin_5026 = frame (4k)
frame_vm_group_bin_5027 = frame (4k)
frame_vm_group_bin_5028 = frame (4k)
frame_vm_group_bin_5029 = frame (4k)
frame_vm_group_bin_5030 = frame (4k)
frame_vm_group_bin_5031 = frame (4k)
frame_vm_group_bin_5032 = frame (4k)
frame_vm_group_bin_5033 = frame (4k)
frame_vm_group_bin_5034 = frame (4k)
frame_vm_group_bin_5035 = frame (4k)
frame_vm_group_bin_5036 = frame (4k)
frame_vm_group_bin_5037 = frame (4k)
frame_vm_group_bin_5038 = frame (4k)
frame_vm_group_bin_5039 = frame (4k)
frame_vm_group_bin_5040 = frame (4k)
frame_vm_group_bin_5041 = frame (4k)
frame_vm_group_bin_5042 = frame (4k)
frame_vm_group_bin_5043 = frame (4k)
frame_vm_group_bin_5044 = frame (4k)
frame_vm_group_bin_5045 = frame (4k)
frame_vm_group_bin_5046 = frame (4k)
frame_vm_group_bin_5047 = frame (4k)
frame_vm_group_bin_5048 = frame (4k)
frame_vm_group_bin_5049 = frame (4k)
frame_vm_group_bin_5050 = frame (4k)
frame_vm_group_bin_5051 = frame (4k)
frame_vm_group_bin_5052 = frame (4k)
frame_vm_group_bin_5053 = frame (4k)
frame_vm_group_bin_5054 = frame (4k)
frame_vm_group_bin_5055 = frame (4k)
frame_vm_group_bin_5056 = frame (4k)
frame_vm_group_bin_5057 = frame (4k)
frame_vm_group_bin_5058 = frame (4k)
frame_vm_group_bin_5059 = frame (4k)
frame_vm_group_bin_5060 = frame (4k)
frame_vm_group_bin_5061 = frame (4k)
frame_vm_group_bin_5062 = frame (4k)
frame_vm_group_bin_5063 = frame (4k)
frame_vm_group_bin_5064 = frame (4k)
frame_vm_group_bin_5065 = frame (4k)
frame_vm_group_bin_5066 = frame (4k)
frame_vm_group_bin_5067 = frame (4k)
frame_vm_group_bin_5068 = frame (4k)
frame_vm_group_bin_5069 = frame (4k)
frame_vm_group_bin_5070 = frame (4k)
frame_vm_group_bin_5071 = frame (4k)
frame_vm_group_bin_5072 = frame (4k)
frame_vm_group_bin_5073 = frame (4k)
frame_vm_group_bin_5074 = frame (4k)
frame_vm_group_bin_5075 = frame (4k)
frame_vm_group_bin_5076 = frame (4k)
frame_vm_group_bin_5077 = frame (4k)
frame_vm_group_bin_5078 = frame (4k)
frame_vm_group_bin_5079 = frame (4k)
frame_vm_group_bin_5080 = frame (4k)
frame_vm_group_bin_5081 = frame (4k)
frame_vm_group_bin_5082 = frame (4k)
frame_vm_group_bin_5083 = frame (4k)
frame_vm_group_bin_5084 = frame (4k)
frame_vm_group_bin_5085 = frame (4k)
frame_vm_group_bin_5086 = frame (4k)
frame_vm_group_bin_5087 = frame (4k)
frame_vm_group_bin_5088 = frame (4k)
frame_vm_group_bin_5089 = frame (4k)
frame_vm_group_bin_5090 = frame (4k)
frame_vm_group_bin_5091 = frame (4k)
frame_vm_group_bin_5092 = frame (4k)
frame_vm_group_bin_5093 = frame (4k)
frame_vm_group_bin_5094 = frame (4k)
frame_vm_group_bin_5095 = frame (4k)
frame_vm_group_bin_5096 = frame (4k)
frame_vm_group_bin_5097 = frame (4k)
frame_vm_group_bin_5098 = frame (4k)
frame_vm_group_bin_5099 = frame (4k)
frame_vm_group_bin_5100 = frame (4k)
frame_vm_group_bin_5101 = frame (4k)
frame_vm_group_bin_5102 = frame (4k)
frame_vm_group_bin_5103 = frame (4k)
frame_vm_group_bin_5104 = frame (4k)
frame_vm_group_bin_5105 = frame (4k)
frame_vm_group_bin_5106 = frame (4k)
frame_vm_group_bin_5107 = frame (4k)
frame_vm_group_bin_5108 = frame (4k)
frame_vm_group_bin_5109 = frame (4k)
frame_vm_group_bin_5110 = frame (4k)
frame_vm_group_bin_5111 = frame (4k)
frame_vm_group_bin_5112 = frame (4k)
frame_vm_group_bin_5113 = frame (4k)
frame_vm_group_bin_5114 = frame (4k)
frame_vm_group_bin_5115 = frame (4k)
frame_vm_group_bin_5116 = frame (4k)
frame_vm_group_bin_5117 = frame (4k)
frame_vm_group_bin_5118 = frame (4k)
frame_vm_group_bin_5119 = frame (4k)
frame_vm_group_bin_5120 = frame (4k)
frame_vm_group_bin_5121 = frame (4k)
frame_vm_group_bin_5122 = frame (4k)
frame_vm_group_bin_5123 = frame (4k)
frame_vm_group_bin_5124 = frame (4k)
frame_vm_group_bin_5125 = frame (4k)
frame_vm_group_bin_5126 = frame (4k)
frame_vm_group_bin_5127 = frame (4k)
frame_vm_group_bin_5128 = frame (4k)
frame_vm_group_bin_5129 = frame (4k)
frame_vm_group_bin_5130 = frame (4k)
frame_vm_group_bin_5131 = frame (4k)
frame_vm_group_bin_5132 = frame (4k)
frame_vm_group_bin_5133 = frame (4k)
frame_vm_group_bin_5134 = frame (4k)
frame_vm_group_bin_5135 = frame (4k)
frame_vm_group_bin_5136 = frame (4k)
frame_vm_group_bin_5137 = frame (4k)
frame_vm_group_bin_5138 = frame (4k)
frame_vm_group_bin_5139 = frame (4k)
frame_vm_group_bin_5140 = frame (4k)
frame_vm_group_bin_5141 = frame (4k)
frame_vm_group_bin_5142 = frame (4k)
frame_vm_group_bin_5143 = frame (4k)
frame_vm_group_bin_5144 = frame (4k)
frame_vm_group_bin_5145 = frame (4k)
frame_vm_group_bin_5146 = frame (4k)
frame_vm_group_bin_5147 = frame (4k)
frame_vm_group_bin_5148 = frame (4k)
frame_vm_group_bin_5149 = frame (4k)
frame_vm_group_bin_5150 = frame (4k)
frame_vm_group_bin_5151 = frame (4k)
frame_vm_group_bin_5152 = frame (4k)
frame_vm_group_bin_5153 = frame (4k)
frame_vm_group_bin_5154 = frame (4k)
frame_vm_group_bin_5155 = frame (4k)
frame_vm_group_bin_5156 = frame (4k)
frame_vm_group_bin_5157 = frame (4k)
frame_vm_group_bin_5158 = frame (4k)
frame_vm_group_bin_5159 = frame (4k)
frame_vm_group_bin_5160 = frame (4k)
frame_vm_group_bin_5161 = frame (4k)
frame_vm_group_bin_5162 = frame (4k)
frame_vm_group_bin_5163 = frame (4k)
frame_vm_group_bin_5164 = frame (4k)
frame_vm_group_bin_5165 = frame (4k)
frame_vm_group_bin_5166 = frame (4k)
frame_vm_group_bin_5167 = frame (4k)
frame_vm_group_bin_5168 = frame (4k)
frame_vm_group_bin_5169 = frame (4k)
frame_vm_group_bin_5170 = frame (4k)
frame_vm_group_bin_5171 = frame (4k)
frame_vm_group_bin_5172 = frame (4k)
frame_vm_group_bin_5173 = frame (4k)
frame_vm_group_bin_5174 = frame (4k)
frame_vm_group_bin_5175 = frame (4k)
frame_vm_group_bin_5176 = frame (4k)
frame_vm_group_bin_5177 = frame (4k)
frame_vm_group_bin_5178 = frame (4k)
frame_vm_group_bin_5179 = frame (4k)
frame_vm_group_bin_5180 = frame (4k)
frame_vm_group_bin_5181 = frame (4k)
frame_vm_group_bin_5182 = frame (4k)
frame_vm_group_bin_5183 = frame (4k)
frame_vm_group_bin_5184 = frame (4k)
frame_vm_group_bin_5185 = frame (4k)
frame_vm_group_bin_5186 = frame (4k)
frame_vm_group_bin_5187 = frame (4k)
frame_vm_group_bin_5188 = frame (4k)
frame_vm_group_bin_5189 = frame (4k)
frame_vm_group_bin_5190 = frame (4k)
frame_vm_group_bin_5191 = frame (4k)
frame_vm_group_bin_5192 = frame (4k)
frame_vm_group_bin_5193 = frame (4k)
frame_vm_group_bin_5194 = frame (4k)
frame_vm_group_bin_5195 = frame (4k)
frame_vm_group_bin_5196 = frame (4k)
frame_vm_group_bin_5197 = frame (4k)
frame_vm_group_bin_5198 = frame (4k)
frame_vm_group_bin_5199 = frame (4k)
frame_vm_group_bin_5200 = frame (4k)
frame_vm_group_bin_5201 = frame (4k)
frame_vm_group_bin_5202 = frame (4k)
frame_vm_group_bin_5203 = frame (4k)
frame_vm_group_bin_5204 = frame (4k)
frame_vm_group_bin_5205 = frame (4k)
frame_vm_group_bin_5206 = frame (4k)
frame_vm_group_bin_5207 = frame (4k)
frame_vm_group_bin_5208 = frame (4k)
frame_vm_group_bin_5209 = frame (4k)
frame_vm_group_bin_5210 = frame (4k)
frame_vm_group_bin_5211 = frame (4k)
frame_vm_group_bin_5212 = frame (4k)
frame_vm_group_bin_5213 = frame (4k)
frame_vm_group_bin_5214 = frame (4k)
frame_vm_group_bin_5215 = frame (4k)
frame_vm_group_bin_5216 = frame (4k)
frame_vm_group_bin_5217 = frame (4k)
frame_vm_group_bin_5218 = frame (4k)
frame_vm_group_bin_5219 = frame (4k)
frame_vm_group_bin_5220 = frame (4k)
frame_vm_group_bin_5221 = frame (4k)
frame_vm_group_bin_5222 = frame (4k)
frame_vm_group_bin_5223 = frame (4k)
frame_vm_group_bin_5224 = frame (4k)
frame_vm_group_bin_5225 = frame (4k)
frame_vm_group_bin_5226 = frame (4k)
frame_vm_group_bin_5227 = frame (4k)
frame_vm_group_bin_5228 = frame (4k)
frame_vm_group_bin_5229 = frame (4k)
frame_vm_group_bin_5230 = frame (4k)
frame_vm_group_bin_5231 = frame (4k)
frame_vm_group_bin_5232 = frame (4k)
frame_vm_group_bin_5233 = frame (4k)
frame_vm_group_bin_5234 = frame (4k)
frame_vm_group_bin_5235 = frame (4k)
frame_vm_group_bin_5236 = frame (4k)
frame_vm_group_bin_5237 = frame (4k)
frame_vm_group_bin_5238 = frame (4k)
frame_vm_group_bin_5239 = frame (4k)
frame_vm_group_bin_5240 = frame (4k)
frame_vm_group_bin_5241 = frame (4k)
frame_vm_group_bin_5242 = frame (4k)
frame_vm_group_bin_5243 = frame (4k)
frame_vm_group_bin_5244 = frame (4k)
frame_vm_group_bin_5245 = frame (4k)
frame_vm_group_bin_5246 = frame (4k)
frame_vm_group_bin_5247 = frame (4k)
frame_vm_group_bin_5248 = frame (4k)
frame_vm_group_bin_5249 = frame (4k)
frame_vm_group_bin_5250 = frame (4k)
frame_vm_group_bin_5251 = frame (4k)
frame_vm_group_bin_5252 = frame (4k)
frame_vm_group_bin_5253 = frame (4k)
frame_vm_group_bin_5254 = frame (4k)
frame_vm_group_bin_5255 = frame (4k)
frame_vm_group_bin_5256 = frame (4k)
frame_vm_group_bin_5257 = frame (4k)
frame_vm_group_bin_5258 = frame (4k)
frame_vm_group_bin_5259 = frame (4k)
frame_vm_group_bin_5260 = frame (4k)
frame_vm_group_bin_5261 = frame (4k)
frame_vm_group_bin_5262 = frame (4k)
frame_vm_group_bin_5263 = frame (4k)
frame_vm_group_bin_5264 = frame (4k)
frame_vm_group_bin_5265 = frame (4k)
frame_vm_group_bin_5266 = frame (4k)
frame_vm_group_bin_5267 = frame (4k)
frame_vm_group_bin_5268 = frame (4k)
frame_vm_group_bin_5269 = frame (4k)
frame_vm_group_bin_5270 = frame (4k)
frame_vm_group_bin_5271 = frame (4k)
frame_vm_group_bin_5272 = frame (4k)
frame_vm_group_bin_5273 = frame (4k)
frame_vm_group_bin_5274 = frame (4k)
frame_vm_group_bin_5275 = frame (4k)
frame_vm_group_bin_5276 = frame (4k)
frame_vm_group_bin_5277 = frame (4k)
frame_vm_group_bin_5278 = frame (4k)
frame_vm_group_bin_5279 = frame (4k)
frame_vm_group_bin_5280 = frame (4k)
frame_vm_group_bin_5281 = frame (4k)
frame_vm_group_bin_5282 = frame (4k)
frame_vm_group_bin_5283 = frame (4k)
frame_vm_group_bin_5284 = frame (4k)
frame_vm_group_bin_5285 = frame (4k)
frame_vm_group_bin_5286 = frame (4k)
frame_vm_group_bin_5287 = frame (4k)
frame_vm_group_bin_5288 = frame (4k)
frame_vm_group_bin_5289 = frame (4k)
frame_vm_group_bin_5290 = frame (4k)
frame_vm_group_bin_5291 = frame (4k)
frame_vm_group_bin_5292 = frame (4k)
frame_vm_group_bin_5293 = frame (4k)
frame_vm_group_bin_5294 = frame (4k)
frame_vm_group_bin_5295 = frame (4k)
frame_vm_group_bin_5297 = frame (4k)
frame_vm_group_bin_5298 = frame (4k)
frame_vm_group_bin_5299 = frame (4k)
frame_vm_group_bin_5300 = frame (4k)
frame_vm_group_bin_5301 = frame (4k)
frame_vm_group_bin_5302 = frame (4k)
frame_vm_group_bin_5303 = frame (4k)
frame_vm_group_bin_5304 = frame (4k)
frame_vm_group_bin_5305 = frame (4k)
frame_vm_group_bin_5306 = frame (4k)
frame_vm_group_bin_5307 = frame (4k)
frame_vm_group_bin_5308 = frame (4k)
frame_vm_group_bin_5309 = frame (4k)
frame_vm_group_bin_5310 = frame (4k)
frame_vm_group_bin_5311 = frame (4k)
frame_vm_group_bin_5312 = frame (4k)
frame_vm_group_bin_5313 = frame (4k)
frame_vm_group_bin_5314 = frame (4k)
frame_vm_group_bin_5315 = frame (4k)
frame_vm_group_bin_5316 = frame (4k)
frame_vm_group_bin_5317 = frame (4k)
frame_vm_group_bin_5318 = frame (4k)
frame_vm_group_bin_5319 = frame (4k)
frame_vm_group_bin_5320 = frame (4k)
frame_vm_group_bin_5321 = frame (4k)
frame_vm_group_bin_5322 = frame (4k)
frame_vm_group_bin_5323 = frame (4k)
frame_vm_group_bin_5324 = frame (4k)
frame_vm_group_bin_5325 = frame (4k)
frame_vm_group_bin_5326 = frame (4k)
frame_vm_group_bin_5327 = frame (4k)
frame_vm_group_bin_5328 = frame (4k)
frame_vm_group_bin_5329 = frame (4k)
frame_vm_group_bin_5330 = frame (4k)
frame_vm_group_bin_5331 = frame (4k)
frame_vm_group_bin_5332 = frame (4k)
frame_vm_group_bin_5333 = frame (4k)
frame_vm_group_bin_5334 = frame (4k)
frame_vm_group_bin_5335 = frame (4k)
frame_vm_group_bin_5336 = frame (4k)
frame_vm_group_bin_5337 = frame (4k)
frame_vm_group_bin_5338 = frame (4k)
frame_vm_group_bin_5339 = frame (4k)
frame_vm_group_bin_5340 = frame (4k)
frame_vm_group_bin_5341 = frame (4k)
frame_vm_group_bin_5342 = frame (4k)
frame_vm_group_bin_5343 = frame (4k)
frame_vm_group_bin_5344 = frame (4k)
frame_vm_group_bin_5345 = frame (4k)
frame_vm_group_bin_5346 = frame (4k)
frame_vm_group_bin_5347 = frame (4k)
frame_vm_group_bin_5348 = frame (4k)
frame_vm_group_bin_5349 = frame (4k)
frame_vm_group_bin_5350 = frame (4k)
frame_vm_group_bin_5351 = frame (4k)
frame_vm_group_bin_5352 = frame (4k)
frame_vm_group_bin_5353 = frame (4k)
frame_vm_group_bin_5354 = frame (4k)
frame_vm_group_bin_5355 = frame (4k)
frame_vm_group_bin_5356 = frame (4k)
frame_vm_group_bin_5357 = frame (4k)
frame_vm_group_bin_5358 = frame (4k)
frame_vm_group_bin_5359 = frame (4k)
frame_vm_group_bin_5360 = frame (4k)
frame_vm_group_bin_5361 = frame (4k)
frame_vm_group_bin_5362 = frame (4k)
frame_vm_group_bin_5363 = frame (4k)
frame_vm_group_bin_5364 = frame (4k)
frame_vm_group_bin_5365 = frame (4k)
frame_vm_group_bin_5366 = frame (4k)
frame_vm_group_bin_5367 = frame (4k)
frame_vm_group_bin_5368 = frame (4k)
frame_vm_group_bin_5369 = frame (4k)
frame_vm_group_bin_5370 = frame (4k)
frame_vm_group_bin_5371 = frame (4k)
frame_vm_group_bin_5372 = frame (4k)
frame_vm_group_bin_5373 = frame (4k)
frame_vm_group_bin_5374 = frame (4k)
frame_vm_group_bin_5375 = frame (4k)
frame_vm_group_bin_5376 = frame (4k)
frame_vm_group_bin_5377 = frame (4k)
frame_vm_group_bin_5378 = frame (4k)
frame_vm_group_bin_5379 = frame (4k)
frame_vm_group_bin_5380 = frame (4k)
frame_vm_group_bin_5381 = frame (4k)
frame_vm_group_bin_5382 = frame (4k)
frame_vm_group_bin_5383 = frame (4k)
frame_vm_group_bin_5384 = frame (4k)
frame_vm_group_bin_5385 = frame (4k)
frame_vm_group_bin_5386 = frame (4k)
frame_vm_group_bin_5387 = frame (4k)
frame_vm_group_bin_5388 = frame (4k)
frame_vm_group_bin_5389 = frame (4k)
frame_vm_group_bin_5390 = frame (4k)
frame_vm_group_bin_5391 = frame (4k)
frame_vm_group_bin_5392 = frame (4k)
frame_vm_group_bin_5393 = frame (4k)
frame_vm_group_bin_5394 = frame (4k)
frame_vm_group_bin_5395 = frame (4k)
frame_vm_group_bin_5396 = frame (4k)
frame_vm_group_bin_5397 = frame (4k)
frame_vm_group_bin_5398 = frame (4k)
frame_vm_group_bin_5399 = frame (4k)
frame_vm_group_bin_5400 = frame (4k)
frame_vm_group_bin_5401 = frame (4k)
frame_vm_group_bin_5402 = frame (4k)
frame_vm_group_bin_5403 = frame (4k)
frame_vm_group_bin_5404 = frame (4k)
frame_vm_group_bin_5405 = frame (4k)
frame_vm_group_bin_5406 = frame (4k)
frame_vm_group_bin_5407 = frame (4k)
frame_vm_group_bin_5408 = frame (4k)
frame_vm_group_bin_5409 = frame (4k)
frame_vm_group_bin_5410 = frame (4k)
frame_vm_group_bin_5411 = frame (4k)
frame_vm_group_bin_5412 = frame (4k)
frame_vm_group_bin_5413 = frame (4k)
frame_vm_group_bin_5414 = frame (4k)
frame_vm_group_bin_5415 = frame (4k)
frame_vm_group_bin_5416 = frame (4k)
frame_vm_group_bin_5417 = frame (4k)
frame_vm_group_bin_5418 = frame (4k)
frame_vm_group_bin_5419 = frame (4k)
frame_vm_group_bin_5420 = frame (4k)
frame_vm_group_bin_5421 = frame (4k)
frame_vm_group_bin_5422 = frame (4k)
frame_vm_group_bin_5423 = frame (4k)
frame_vm_group_bin_5424 = frame (4k)
frame_vm_group_bin_5425 = frame (4k)
frame_vm_group_bin_5426 = frame (4k)
frame_vm_group_bin_5427 = frame (4k)
frame_vm_group_bin_5428 = frame (4k)
frame_vm_group_bin_5429 = frame (4k)
frame_vm_group_bin_5430 = frame (4k)
frame_vm_group_bin_5431 = frame (4k)
frame_vm_group_bin_5432 = frame (4k)
frame_vm_group_bin_5433 = frame (4k)
frame_vm_group_bin_5434 = frame (4k)
frame_vm_group_bin_5435 = frame (4k)
frame_vm_group_bin_5436 = frame (4k)
frame_vm_group_bin_5437 = frame (4k)
frame_vm_group_bin_5438 = frame (4k)
frame_vm_group_bin_5439 = frame (4k)
frame_vm_group_bin_5440 = frame (4k)
frame_vm_group_bin_5441 = frame (4k)
frame_vm_group_bin_5442 = frame (4k)
frame_vm_group_bin_5443 = frame (4k)
frame_vm_group_bin_5444 = frame (4k)
frame_vm_group_bin_5445 = frame (4k)
frame_vm_group_bin_5446 = frame (4k)
frame_vm_group_bin_5447 = frame (4k)
frame_vm_group_bin_5448 = frame (4k)
frame_vm_group_bin_5449 = frame (4k)
frame_vm_group_bin_5450 = frame (4k)
frame_vm_group_bin_5451 = frame (4k)
frame_vm_group_bin_5452 = frame (4k)
frame_vm_group_bin_5453 = frame (4k)
frame_vm_group_bin_5454 = frame (4k)
frame_vm_group_bin_5455 = frame (4k)
frame_vm_group_bin_5456 = frame (4k)
frame_vm_group_bin_5457 = frame (4k)
frame_vm_group_bin_5458 = frame (4k)
frame_vm_group_bin_5459 = frame (4k)
frame_vm_group_bin_5460 = frame (4k)
frame_vm_group_bin_5461 = frame (4k)
frame_vm_group_bin_5462 = frame (4k)
frame_vm_group_bin_5463 = frame (4k)
frame_vm_group_bin_5464 = frame (4k)
frame_vm_group_bin_5465 = frame (4k)
frame_vm_group_bin_5466 = frame (4k)
frame_vm_group_bin_5467 = frame (4k)
frame_vm_group_bin_5468 = frame (4k)
frame_vm_group_bin_5469 = frame (4k)
frame_vm_group_bin_5470 = frame (4k)
frame_vm_group_bin_5471 = frame (4k)
frame_vm_group_bin_5472 = frame (4k)
frame_vm_group_bin_5473 = frame (4k)
frame_vm_group_bin_5474 = frame (4k)
frame_vm_group_bin_5475 = frame (4k)
frame_vm_group_bin_5476 = frame (4k)
frame_vm_group_bin_5477 = frame (4k)
frame_vm_group_bin_5478 = frame (4k)
frame_vm_group_bin_5479 = frame (4k)
frame_vm_group_bin_5480 = frame (4k)
frame_vm_group_bin_5481 = frame (4k)
frame_vm_group_bin_5482 = frame (4k)
frame_vm_group_bin_5483 = frame (4k)
frame_vm_group_bin_5484 = frame (4k)
frame_vm_group_bin_5485 = frame (4k)
frame_vm_group_bin_5486 = frame (4k)
frame_vm_group_bin_5487 = frame (4k)
frame_vm_group_bin_5488 = frame (4k)
frame_vm_group_bin_5489 = frame (4k)
frame_vm_group_bin_5490 = frame (4k)
frame_vm_group_bin_5491 = frame (4k)
frame_vm_group_bin_5492 = frame (4k)
frame_vm_group_bin_5493 = frame (4k)
frame_vm_group_bin_5494 = frame (4k)
frame_vm_group_bin_5495 = frame (4k)
frame_vm_group_bin_5496 = frame (4k)
frame_vm_group_bin_5497 = frame (4k)
frame_vm_group_bin_5498 = frame (4k)
frame_vm_group_bin_5499 = frame (4k)
frame_vm_group_bin_5500 = frame (4k)
frame_vm_group_bin_5501 = frame (4k)
frame_vm_group_bin_5502 = frame (4k)
frame_vm_group_bin_5503 = frame (4k)
frame_vm_group_bin_5504 = frame (4k)
frame_vm_group_bin_5505 = frame (4k)
frame_vm_group_bin_5506 = frame (4k)
frame_vm_group_bin_5507 = frame (4k)
frame_vm_group_bin_5508 = frame (4k)
frame_vm_group_bin_5509 = frame (4k)
frame_vm_group_bin_5510 = frame (4k)
frame_vm_group_bin_5511 = frame (4k)
frame_vm_group_bin_5512 = frame (4k)
frame_vm_group_bin_5513 = frame (4k)
frame_vm_group_bin_5514 = frame (4k)
frame_vm_group_bin_5515 = frame (4k)
frame_vm_group_bin_5516 = frame (4k)
frame_vm_group_bin_5517 = frame (4k)
frame_vm_group_bin_5518 = frame (4k)
frame_vm_group_bin_5519 = frame (4k)
frame_vm_group_bin_5520 = frame (4k)
frame_vm_group_bin_5521 = frame (4k)
frame_vm_group_bin_5522 = frame (4k)
frame_vm_group_bin_5523 = frame (4k)
frame_vm_group_bin_5524 = frame (4k)
frame_vm_group_bin_5525 = frame (4k)
frame_vm_group_bin_5526 = frame (4k)
frame_vm_group_bin_5527 = frame (4k)
frame_vm_group_bin_5528 = frame (4k)
frame_vm_group_bin_5529 = frame (4k)
frame_vm_group_bin_5530 = frame (4k)
frame_vm_group_bin_5531 = frame (4k)
frame_vm_group_bin_5532 = frame (4k)
frame_vm_group_bin_5533 = frame (4k)
frame_vm_group_bin_5534 = frame (4k)
frame_vm_group_bin_5535 = frame (4k)
frame_vm_group_bin_5536 = frame (4k)
frame_vm_group_bin_5537 = frame (4k)
frame_vm_group_bin_5538 = frame (4k)
frame_vm_group_bin_5539 = frame (4k)
frame_vm_group_bin_5540 = frame (4k)
frame_vm_group_bin_5541 = frame (4k)
frame_vm_group_bin_5542 = frame (4k)
frame_vm_group_bin_5543 = frame (4k)
frame_vm_group_bin_5544 = frame (4k)
frame_vm_group_bin_5545 = frame (4k)
frame_vm_group_bin_5546 = frame (4k)
frame_vm_group_bin_5547 = frame (4k)
frame_vm_group_bin_5548 = frame (4k)
frame_vm_group_bin_5549 = frame (4k)
frame_vm_group_bin_5550 = frame (4k)
frame_vm_group_bin_5551 = frame (4k)
frame_vm_group_bin_5552 = frame (4k)
frame_vm_group_bin_5553 = frame (4k)
frame_vm_group_bin_5554 = frame (4k)
frame_vm_group_bin_5555 = frame (4k)
frame_vm_group_bin_5556 = frame (4k)
frame_vm_group_bin_5557 = frame (4k)
frame_vm_group_bin_5558 = frame (4k)
frame_vm_group_bin_5559 = frame (4k)
frame_vm_group_bin_5560 = frame (4k)
frame_vm_group_bin_5561 = frame (4k)
frame_vm_group_bin_5562 = frame (4k)
frame_vm_group_bin_5563 = frame (4k)
frame_vm_group_bin_5564 = frame (4k)
frame_vm_group_bin_5565 = frame (4k)
frame_vm_group_bin_5566 = frame (4k)
frame_vm_group_bin_5567 = frame (4k)
frame_vm_group_bin_5568 = frame (4k)
frame_vm_group_bin_5569 = frame (4k)
frame_vm_group_bin_5570 = frame (4k)
frame_vm_group_bin_5571 = frame (4k)
frame_vm_group_bin_5572 = frame (4k)
frame_vm_group_bin_5573 = frame (4k)
frame_vm_group_bin_5574 = frame (4k)
frame_vm_group_bin_5575 = frame (4k)
frame_vm_group_bin_5576 = frame (4k)
frame_vm_group_bin_5577 = frame (4k)
frame_vm_group_bin_5578 = frame (4k)
frame_vm_group_bin_5579 = frame (4k)
frame_vm_group_bin_5580 = frame (4k)
frame_vm_group_bin_5581 = frame (4k)
frame_vm_group_bin_5582 = frame (4k)
frame_vm_group_bin_5583 = frame (4k)
frame_vm_group_bin_5584 = frame (4k)
frame_vm_group_bin_5585 = frame (4k)
frame_vm_group_bin_5586 = frame (4k)
frame_vm_group_bin_5587 = frame (4k)
frame_vm_group_bin_5588 = frame (4k)
frame_vm_group_bin_5589 = frame (4k)
frame_vm_group_bin_5590 = frame (4k)
frame_vm_group_bin_5591 = frame (4k)
frame_vm_group_bin_5592 = frame (4k)
frame_vm_group_bin_5593 = frame (4k)
frame_vm_group_bin_5594 = frame (4k)
frame_vm_group_bin_5595 = frame (4k)
frame_vm_group_bin_5596 = frame (4k)
frame_vm_group_bin_5597 = frame (4k)
frame_vm_group_bin_5598 = frame (4k)
frame_vm_group_bin_5599 = frame (4k)
frame_vm_group_bin_5600 = frame (4k)
frame_vm_group_bin_5601 = frame (4k)
frame_vm_group_bin_5602 = frame (4k)
frame_vm_group_bin_5603 = frame (4k)
frame_vm_group_bin_5604 = frame (4k)
frame_vm_group_bin_5605 = frame (4k)
frame_vm_group_bin_5606 = frame (4k)
frame_vm_group_bin_5607 = frame (4k)
frame_vm_group_bin_5608 = frame (4k)
frame_vm_group_bin_5609 = frame (4k)
frame_vm_group_bin_5610 = frame (4k)
frame_vm_group_bin_5611 = frame (4k)
frame_vm_group_bin_5612 = frame (4k)
frame_vm_group_bin_5613 = frame (4k)
frame_vm_group_bin_5614 = frame (4k)
frame_vm_group_bin_5615 = frame (4k)
frame_vm_group_bin_5616 = frame (4k)
frame_vm_group_bin_5617 = frame (4k)
frame_vm_group_bin_5618 = frame (4k)
frame_vm_group_bin_5619 = frame (4k)
frame_vm_group_bin_5620 = frame (4k)
frame_vm_group_bin_5621 = frame (4k)
frame_vm_group_bin_5622 = frame (4k)
frame_vm_group_bin_5623 = frame (4k)
frame_vm_group_bin_5624 = frame (4k)
frame_vm_group_bin_5625 = frame (4k)
frame_vm_group_bin_5626 = frame (4k)
frame_vm_group_bin_5627 = frame (4k)
frame_vm_group_bin_5628 = frame (4k)
frame_vm_group_bin_5629 = frame (4k)
frame_vm_group_bin_5630 = frame (4k)
frame_vm_group_bin_5631 = frame (4k)
frame_vm_group_bin_5632 = frame (4k)
frame_vm_group_bin_5633 = frame (4k)
frame_vm_group_bin_5634 = frame (4k)
frame_vm_group_bin_5635 = frame (4k)
frame_vm_group_bin_5636 = frame (4k)
frame_vm_group_bin_5637 = frame (4k)
frame_vm_group_bin_5638 = frame (4k)
frame_vm_group_bin_5639 = frame (4k)
frame_vm_group_bin_5640 = frame (4k)
frame_vm_group_bin_5641 = frame (4k)
frame_vm_group_bin_5642 = frame (4k)
frame_vm_group_bin_5643 = frame (4k)
frame_vm_group_bin_5644 = frame (4k)
frame_vm_group_bin_5645 = frame (4k)
frame_vm_group_bin_5646 = frame (4k)
frame_vm_group_bin_5647 = frame (4k)
frame_vm_group_bin_5648 = frame (4k)
frame_vm_group_bin_5649 = frame (4k)
frame_vm_group_bin_5650 = frame (4k)
frame_vm_group_bin_5651 = frame (4k)
frame_vm_group_bin_5652 = frame (4k)
frame_vm_group_bin_5653 = frame (4k)
frame_vm_group_bin_5654 = frame (4k)
frame_vm_group_bin_5655 = frame (4k)
frame_vm_group_bin_5656 = frame (4k)
frame_vm_group_bin_5657 = frame (4k)
frame_vm_group_bin_5658 = frame (4k)
frame_vm_group_bin_5659 = frame (4k)
frame_vm_group_bin_5660 = frame (4k)
frame_vm_group_bin_5661 = frame (4k)
frame_vm_group_bin_5662 = frame (4k)
frame_vm_group_bin_5663 = frame (4k)
frame_vm_group_bin_5664 = frame (4k)
frame_vm_group_bin_5665 = frame (4k)
frame_vm_group_bin_5666 = frame (4k)
frame_vm_group_bin_5667 = frame (4k)
frame_vm_group_bin_5668 = frame (4k)
frame_vm_group_bin_5669 = frame (4k)
frame_vm_group_bin_5670 = frame (4k)
frame_vm_group_bin_5671 = frame (4k)
frame_vm_group_bin_5672 = frame (4k)
frame_vm_group_bin_5673 = frame (4k)
frame_vm_group_bin_5674 = frame (4k)
frame_vm_group_bin_5675 = frame (4k)
frame_vm_group_bin_5676 = frame (4k)
frame_vm_group_bin_5677 = frame (4k)
frame_vm_group_bin_5678 = frame (4k)
frame_vm_group_bin_5679 = frame (4k)
frame_vm_group_bin_5680 = frame (4k)
frame_vm_group_bin_5681 = frame (4k)
frame_vm_group_bin_5682 = frame (4k)
frame_vm_group_bin_5683 = frame (4k)
frame_vm_group_bin_5684 = frame (4k)
frame_vm_group_bin_5685 = frame (4k)
frame_vm_group_bin_5686 = frame (4k)
frame_vm_group_bin_5687 = frame (4k)
frame_vm_group_bin_5688 = frame (4k)
frame_vm_group_bin_5689 = frame (4k)
frame_vm_group_bin_5690 = frame (4k)
frame_vm_group_bin_5691 = frame (4k)
frame_vm_group_bin_5692 = frame (4k)
frame_vm_group_bin_5693 = frame (4k)
frame_vm_group_bin_5694 = frame (4k)
frame_vm_group_bin_5695 = frame (4k)
frame_vm_group_bin_5696 = frame (4k)
frame_vm_group_bin_5697 = frame (4k)
frame_vm_group_bin_5698 = frame (4k)
frame_vm_group_bin_5699 = frame (4k)
frame_vm_group_bin_5700 = frame (4k)
frame_vm_group_bin_5701 = frame (4k)
frame_vm_group_bin_5702 = frame (4k)
frame_vm_group_bin_5703 = frame (4k)
frame_vm_group_bin_5704 = frame (4k)
frame_vm_group_bin_5705 = frame (4k)
frame_vm_group_bin_5706 = frame (4k)
frame_vm_group_bin_5707 = frame (4k)
frame_vm_group_bin_5708 = frame (4k)
frame_vm_group_bin_5709 = frame (4k)
frame_vm_group_bin_5710 = frame (4k)
frame_vm_group_bin_5711 = frame (4k)
frame_vm_group_bin_5712 = frame (4k)
frame_vm_group_bin_5713 = frame (4k)
frame_vm_group_bin_5714 = frame (4k)
frame_vm_group_bin_5715 = frame (4k)
frame_vm_group_bin_5716 = frame (4k)
frame_vm_group_bin_5717 = frame (4k)
frame_vm_group_bin_5718 = frame (4k)
frame_vm_group_bin_5719 = frame (4k)
frame_vm_group_bin_5720 = frame (4k)
frame_vm_group_bin_5721 = frame (4k)
frame_vm_group_bin_5722 = frame (4k)
frame_vm_group_bin_5723 = frame (4k)
frame_vm_group_bin_5724 = frame (4k)
frame_vm_group_bin_5725 = frame (4k)
frame_vm_group_bin_5726 = frame (4k)
frame_vm_group_bin_5727 = frame (4k)
frame_vm_group_bin_5728 = frame (4k)
frame_vm_group_bin_5729 = frame (4k)
frame_vm_group_bin_5730 = frame (4k)
frame_vm_group_bin_5731 = frame (4k)
frame_vm_group_bin_5732 = frame (4k)
frame_vm_group_bin_5733 = frame (4k)
frame_vm_group_bin_5734 = frame (4k)
frame_vm_group_bin_5735 = frame (4k)
frame_vm_group_bin_5736 = frame (4k)
frame_vm_group_bin_5737 = frame (4k)
frame_vm_group_bin_5738 = frame (4k)
frame_vm_group_bin_5739 = frame (4k)
frame_vm_group_bin_5740 = frame (4k)
frame_vm_group_bin_5741 = frame (4k)
frame_vm_group_bin_5742 = frame (4k)
frame_vm_group_bin_5743 = frame (4k)
frame_vm_group_bin_5744 = frame (4k)
frame_vm_group_bin_5745 = frame (4k)
frame_vm_group_bin_5746 = frame (4k)
frame_vm_group_bin_5747 = frame (4k)
frame_vm_group_bin_5748 = frame (4k)
frame_vm_group_bin_5749 = frame (4k)
frame_vm_group_bin_5750 = frame (4k)
frame_vm_group_bin_5751 = frame (4k)
frame_vm_group_bin_5752 = frame (4k)
frame_vm_group_bin_5753 = frame (4k)
frame_vm_group_bin_5754 = frame (4k)
frame_vm_group_bin_5755 = frame (4k)
frame_vm_group_bin_5756 = frame (4k)
frame_vm_group_bin_5757 = frame (4k)
frame_vm_group_bin_5758 = frame (4k)
frame_vm_group_bin_5759 = frame (4k)
frame_vm_group_bin_5760 = frame (4k)
frame_vm_group_bin_5761 = frame (4k)
frame_vm_group_bin_5762 = frame (4k)
frame_vm_group_bin_5763 = frame (4k)
frame_vm_group_bin_5764 = frame (4k)
frame_vm_group_bin_5765 = frame (4k)
frame_vm_group_bin_5766 = frame (4k)
frame_vm_group_bin_5767 = frame (4k)
frame_vm_group_bin_5768 = frame (4k)
frame_vm_group_bin_5769 = frame (4k)
frame_vm_group_bin_5770 = frame (4k)
frame_vm_group_bin_5771 = frame (4k)
frame_vm_group_bin_5772 = frame (4k)
frame_vm_group_bin_5773 = frame (4k)
frame_vm_group_bin_5774 = frame (4k)
frame_vm_group_bin_5775 = frame (4k)
frame_vm_group_bin_5776 = frame (4k)
frame_vm_group_bin_5777 = frame (4k)
frame_vm_group_bin_5778 = frame (4k)
frame_vm_group_bin_5779 = frame (4k)
frame_vm_group_bin_5780 = frame (4k)
frame_vm_group_bin_5781 = frame (4k)
frame_vm_group_bin_5782 = frame (4k)
frame_vm_group_bin_5783 = frame (4k)
frame_vm_group_bin_5784 = frame (4k)
frame_vm_group_bin_5785 = frame (4k)
frame_vm_group_bin_5786 = frame (4k)
frame_vm_group_bin_5787 = frame (4k)
frame_vm_group_bin_5788 = frame (4k)
frame_vm_group_bin_5789 = frame (4k)
frame_vm_group_bin_5790 = frame (4k)
frame_vm_group_bin_5791 = frame (4k)
frame_vm_group_bin_5792 = frame (4k)
frame_vm_group_bin_5793 = frame (4k)
frame_vm_group_bin_5794 = frame (4k)
frame_vm_group_bin_5795 = frame (4k)
frame_vm_group_bin_5796 = frame (4k)
frame_vm_group_bin_5797 = frame (4k)
frame_vm_group_bin_5798 = frame (4k)
frame_vm_group_bin_5799 = frame (4k)
frame_vm_group_bin_5800 = frame (4k)
frame_vm_group_bin_5801 = frame (4k)
frame_vm_group_bin_5802 = frame (4k)
frame_vm_group_bin_5803 = frame (4k)
frame_vm_group_bin_5804 = frame (4k)
frame_vm_group_bin_5805 = frame (4k)
frame_vm_group_bin_5806 = frame (4k)
frame_vm_group_bin_5807 = frame (4k)
frame_vm_group_bin_5808 = frame (4k)
frame_vm_group_bin_5809 = frame (4k)
frame_vm_group_bin_5810 = frame (4k)
frame_vm_group_bin_5811 = frame (4k)
frame_vm_group_bin_5812 = frame (4k)
frame_vm_group_bin_5813 = frame (4k)
frame_vm_group_bin_5814 = frame (4k)
frame_vm_group_bin_5815 = frame (4k)
frame_vm_group_bin_5816 = frame (4k)
frame_vm_group_bin_5817 = frame (4k)
frame_vm_group_bin_5818 = frame (4k)
frame_vm_group_bin_5819 = frame (4k)
frame_vm_group_bin_5820 = frame (4k)
frame_vm_group_bin_5821 = frame (4k)
frame_vm_group_bin_5822 = frame (4k)
frame_vm_group_bin_5823 = frame (4k)
frame_vm_group_bin_5824 = frame (4k)
frame_vm_group_bin_5825 = frame (4k)
frame_vm_group_bin_5826 = frame (4k)
frame_vm_group_bin_5827 = frame (4k)
frame_vm_group_bin_5828 = frame (4k)
frame_vm_group_bin_5829 = frame (4k)
frame_vm_group_bin_5830 = frame (4k)
frame_vm_group_bin_5831 = frame (4k)
frame_vm_group_bin_5832 = frame (4k)
frame_vm_group_bin_5833 = frame (4k)
frame_vm_group_bin_5834 = frame (4k)
frame_vm_group_bin_5835 = frame (4k)
frame_vm_group_bin_5836 = frame (4k)
frame_vm_group_bin_5837 = frame (4k)
frame_vm_group_bin_5838 = frame (4k)
frame_vm_group_bin_5839 = frame (4k)
frame_vm_group_bin_5840 = frame (4k)
frame_vm_group_bin_5841 = frame (4k)
frame_vm_group_bin_5842 = frame (4k)
frame_vm_group_bin_5843 = frame (4k)
frame_vm_group_bin_5844 = frame (4k)
frame_vm_group_bin_5845 = frame (4k)
frame_vm_group_bin_5846 = frame (4k)
frame_vm_group_bin_5847 = frame (4k)
frame_vm_group_bin_5848 = frame (4k)
frame_vm_group_bin_5849 = frame (4k)
frame_vm_group_bin_5850 = frame (4k)
frame_vm_group_bin_5851 = frame (4k)
frame_vm_group_bin_5852 = frame (4k)
frame_vm_group_bin_5853 = frame (4k)
frame_vm_group_bin_5854 = frame (4k)
frame_vm_group_bin_5855 = frame (4k)
frame_vm_group_bin_5856 = frame (4k)
frame_vm_group_bin_5857 = frame (4k)
frame_vm_group_bin_5858 = frame (4k)
frame_vm_group_bin_5859 = frame (4k)
frame_vm_group_bin_5860 = frame (4k)
frame_vm_group_bin_5861 = frame (4k)
frame_vm_group_bin_5862 = frame (4k)
frame_vm_group_bin_5863 = frame (4k)
frame_vm_group_bin_5864 = frame (4k)
frame_vm_group_bin_5865 = frame (4k)
frame_vm_group_bin_5866 = frame (4k)
frame_vm_group_bin_5867 = frame (4k)
frame_vm_group_bin_5868 = frame (4k)
frame_vm_group_bin_5869 = frame (4k)
frame_vm_group_bin_5870 = frame (4k)
frame_vm_group_bin_5871 = frame (4k)
frame_vm_group_bin_5872 = frame (4k)
frame_vm_group_bin_5873 = frame (4k)
frame_vm_group_bin_5874 = frame (4k)
frame_vm_group_bin_5875 = frame (4k)
frame_vm_group_bin_5876 = frame (4k)
frame_vm_group_bin_5877 = frame (4k)
frame_vm_group_bin_5878 = frame (4k)
frame_vm_group_bin_5879 = frame (4k)
frame_vm_group_bin_5880 = frame (4k)
frame_vm_group_bin_5881 = frame (4k)
frame_vm_group_bin_5882 = frame (4k)
frame_vm_group_bin_5883 = frame (4k)
frame_vm_group_bin_5884 = frame (4k)
frame_vm_group_bin_5885 = frame (4k)
frame_vm_group_bin_5886 = frame (4k)
frame_vm_group_bin_5887 = frame (4k)
frame_vm_group_bin_5888 = frame (4k)
frame_vm_group_bin_5889 = frame (4k)
frame_vm_group_bin_5890 = frame (4k)
frame_vm_group_bin_5891 = frame (4k)
frame_vm_group_bin_5892 = frame (4k)
frame_vm_group_bin_5893 = frame (4k)
frame_vm_group_bin_5894 = frame (4k)
frame_vm_group_bin_5895 = frame (4k)
frame_vm_group_bin_5896 = frame (4k)
frame_vm_group_bin_5897 = frame (4k)
frame_vm_group_bin_5898 = frame (4k)
frame_vm_group_bin_5899 = frame (4k)
frame_vm_group_bin_5900 = frame (4k)
frame_vm_group_bin_5901 = frame (4k)
frame_vm_group_bin_5902 = frame (4k)
frame_vm_group_bin_5903 = frame (4k)
frame_vm_group_bin_5904 = frame (4k)
frame_vm_group_bin_5905 = frame (4k)
frame_vm_group_bin_5906 = frame (4k)
frame_vm_group_bin_5907 = frame (4k)
frame_vm_group_bin_5908 = frame (4k)
frame_vm_group_bin_5909 = frame (4k)
frame_vm_group_bin_5910 = frame (4k)
frame_vm_group_bin_5911 = frame (4k)
frame_vm_group_bin_5912 = frame (4k)
frame_vm_group_bin_5913 = frame (4k)
frame_vm_group_bin_5914 = frame (4k)
frame_vm_group_bin_5915 = frame (4k)
frame_vm_group_bin_5916 = frame (4k)
frame_vm_group_bin_5917 = frame (4k)
frame_vm_group_bin_5918 = frame (4k)
frame_vm_group_bin_5919 = frame (4k)
frame_vm_group_bin_5920 = frame (4k)
frame_vm_group_bin_5921 = frame (4k)
frame_vm_group_bin_5922 = frame (4k)
frame_vm_group_bin_5923 = frame (4k)
frame_vm_group_bin_5924 = frame (4k)
frame_vm_group_bin_5925 = frame (4k)
frame_vm_group_bin_5926 = frame (4k)
frame_vm_group_bin_5927 = frame (4k)
frame_vm_group_bin_5928 = frame (4k)
frame_vm_group_bin_5929 = frame (4k)
frame_vm_group_bin_5930 = frame (4k)
frame_vm_group_bin_5931 = frame (4k)
frame_vm_group_bin_5932 = frame (4k)
frame_vm_group_bin_5933 = frame (4k)
frame_vm_group_bin_5934 = frame (4k)
frame_vm_group_bin_5935 = frame (4k)
frame_vm_group_bin_5936 = frame (4k)
frame_vm_group_bin_5937 = frame (4k)
frame_vm_group_bin_5938 = frame (4k)
frame_vm_group_bin_5939 = frame (4k)
frame_vm_group_bin_5940 = frame (4k)
frame_vm_group_bin_5941 = frame (4k)
frame_vm_group_bin_5942 = frame (4k)
frame_vm_group_bin_5943 = frame (4k)
frame_vm_group_bin_5944 = frame (4k)
frame_vm_group_bin_5945 = frame (4k)
frame_vm_group_bin_5946 = frame (4k)
frame_vm_group_bin_5947 = frame (4k)
frame_vm_group_bin_5948 = frame (4k)
frame_vm_group_bin_5949 = frame (4k)
frame_vm_group_bin_5950 = frame (4k)
frame_vm_group_bin_5951 = frame (4k)
frame_vm_group_bin_5952 = frame (4k)
frame_vm_group_bin_5953 = frame (4k)
frame_vm_group_bin_5954 = frame (4k)
frame_vm_group_bin_5955 = frame (4k)
frame_vm_group_bin_5956 = frame (4k)
frame_vm_group_bin_5957 = frame (4k)
frame_vm_group_bin_5958 = frame (4k)
frame_vm_group_bin_5959 = frame (4k)
frame_vm_group_bin_5960 = frame (4k)
frame_vm_group_bin_5961 = frame (4k)
frame_vm_group_bin_5962 = frame (4k)
frame_vm_group_bin_5963 = frame (4k)
frame_vm_group_bin_5964 = frame (4k)
frame_vm_group_bin_5965 = frame (4k)
frame_vm_group_bin_5966 = frame (4k)
frame_vm_group_bin_5967 = frame (4k)
frame_vm_group_bin_5968 = frame (4k)
frame_vm_group_bin_5969 = frame (4k)
frame_vm_group_bin_5970 = frame (4k)
frame_vm_group_bin_5971 = frame (4k)
frame_vm_group_bin_5972 = frame (4k)
frame_vm_group_bin_5973 = frame (4k)
frame_vm_group_bin_5974 = frame (4k)
frame_vm_group_bin_5975 = frame (4k)
frame_vm_group_bin_5976 = frame (4k)
frame_vm_group_bin_5977 = frame (4k)
frame_vm_group_bin_5978 = frame (4k)
frame_vm_group_bin_5979 = frame (4k)
frame_vm_group_bin_5980 = frame (4k)
frame_vm_group_bin_5981 = frame (4k)
frame_vm_group_bin_5982 = frame (4k)
frame_vm_group_bin_5983 = frame (4k)
frame_vm_group_bin_5984 = frame (4k)
frame_vm_group_bin_5985 = frame (4k)
frame_vm_group_bin_5986 = frame (4k)
frame_vm_group_bin_5987 = frame (4k)
frame_vm_group_bin_5988 = frame (4k)
frame_vm_group_bin_5989 = frame (4k)
frame_vm_group_bin_5990 = frame (4k)
frame_vm_group_bin_5991 = frame (4k)
frame_vm_group_bin_5992 = frame (4k)
frame_vm_group_bin_5993 = frame (4k)
frame_vm_group_bin_5994 = frame (4k)
frame_vm_group_bin_5995 = frame (4k)
frame_vm_group_bin_5996 = frame (4k)
frame_vm_group_bin_5997 = frame (4k)
frame_vm_group_bin_5998 = frame (4k)
frame_vm_group_bin_5999 = frame (4k)
frame_vm_group_bin_6000 = frame (4k)
frame_vm_group_bin_6001 = frame (4k)
frame_vm_group_bin_6002 = frame (4k)
frame_vm_group_bin_6003 = frame (4k)
frame_vm_group_bin_6004 = frame (4k)
frame_vm_group_bin_6005 = frame (4k)
frame_vm_group_bin_6006 = frame (4k)
frame_vm_group_bin_6007 = frame (4k)
frame_vm_group_bin_6008 = frame (4k)
frame_vm_group_bin_6009 = frame (4k)
frame_vm_group_bin_6010 = frame (4k)
frame_vm_group_bin_6011 = frame (4k)
frame_vm_group_bin_6012 = frame (4k)
frame_vm_group_bin_6013 = frame (4k)
frame_vm_group_bin_6014 = frame (4k)
frame_vm_group_bin_6015 = frame (4k)
frame_vm_group_bin_6016 = frame (4k)
frame_vm_group_bin_6017 = frame (4k)
frame_vm_group_bin_6018 = frame (4k)
frame_vm_group_bin_6019 = frame (4k)
frame_vm_group_bin_6020 = frame (4k)
frame_vm_group_bin_6021 = frame (4k)
frame_vm_group_bin_6022 = frame (4k)
frame_vm_group_bin_6023 = frame (4k)
frame_vm_group_bin_6024 = frame (4k)
frame_vm_group_bin_6025 = frame (4k)
frame_vm_group_bin_6026 = frame (4k)
frame_vm_group_bin_6027 = frame (4k)
frame_vm_group_bin_6028 = frame (4k)
frame_vm_group_bin_6029 = frame (4k)
frame_vm_group_bin_6030 = frame (4k)
frame_vm_group_bin_6031 = frame (4k)
frame_vm_group_bin_6032 = frame (4k)
frame_vm_group_bin_6033 = frame (4k)
frame_vm_group_bin_6034 = frame (4k)
frame_vm_group_bin_6035 = frame (4k)
frame_vm_group_bin_6036 = frame (4k)
frame_vm_group_bin_6037 = frame (4k)
frame_vm_group_bin_6038 = frame (4k)
frame_vm_group_bin_6039 = frame (4k)
frame_vm_group_bin_6040 = frame (4k)
frame_vm_group_bin_6041 = frame (4k)
frame_vm_group_bin_6042 = frame (4k)
frame_vm_group_bin_6043 = frame (4k)
frame_vm_group_bin_6044 = frame (4k)
frame_vm_group_bin_6045 = frame (4k)
frame_vm_group_bin_6046 = frame (4k)
frame_vm_group_bin_6047 = frame (4k)
frame_vm_group_bin_6048 = frame (4k)
frame_vm_group_bin_6049 = frame (4k)
frame_vm_group_bin_6050 = frame (4k)
frame_vm_group_bin_6051 = frame (4k)
frame_vm_group_bin_6052 = frame (4k)
frame_vm_group_bin_6053 = frame (4k)
frame_vm_group_bin_6054 = frame (4k)
frame_vm_group_bin_6055 = frame (4k)
frame_vm_group_bin_6056 = frame (4k)
frame_vm_group_bin_6057 = frame (4k)
frame_vm_group_bin_6058 = frame (4k)
frame_vm_group_bin_6059 = frame (4k)
frame_vm_group_bin_6060 = frame (4k)
frame_vm_group_bin_6061 = frame (4k)
frame_vm_group_bin_6062 = frame (4k)
frame_vm_group_bin_6063 = frame (4k)
frame_vm_group_bin_6064 = frame (4k)
frame_vm_group_bin_6065 = frame (4k)
frame_vm_group_bin_6066 = frame (4k)
frame_vm_group_bin_6067 = frame (4k)
frame_vm_group_bin_6068 = frame (4k)
frame_vm_group_bin_6069 = frame (4k)
frame_vm_group_bin_6070 = frame (4k)
frame_vm_group_bin_6071 = frame (4k)
frame_vm_group_bin_6072 = frame (4k)
frame_vm_group_bin_6073 = frame (4k)
frame_vm_group_bin_6074 = frame (4k)
frame_vm_group_bin_6075 = frame (4k)
frame_vm_group_bin_6076 = frame (4k)
frame_vm_group_bin_6077 = frame (4k)
frame_vm_group_bin_6078 = frame (4k)
frame_vm_group_bin_6079 = frame (4k)
frame_vm_group_bin_6080 = frame (4k)
frame_vm_group_bin_6081 = frame (4k)
frame_vm_group_bin_6082 = frame (4k)
frame_vm_group_bin_6083 = frame (4k)
frame_vm_group_bin_6084 = frame (4k)
frame_vm_group_bin_6085 = frame (4k)
frame_vm_group_bin_6086 = frame (4k)
frame_vm_group_bin_6087 = frame (4k)
frame_vm_group_bin_6088 = frame (4k)
frame_vm_group_bin_6089 = frame (4k)
frame_vm_group_bin_6090 = frame (4k)
frame_vm_group_bin_6091 = frame (4k)
frame_vm_group_bin_6092 = frame (4k)
frame_vm_group_bin_6093 = frame (4k)
frame_vm_group_bin_6094 = frame (4k)
frame_vm_group_bin_6095 = frame (4k)
frame_vm_group_bin_6096 = frame (4k)
frame_vm_group_bin_6097 = frame (4k)
frame_vm_group_bin_6098 = frame (4k)
frame_vm_group_bin_6099 = frame (4k)
frame_vm_group_bin_6100 = frame (4k)
frame_vm_group_bin_6101 = frame (4k)
frame_vm_group_bin_6102 = frame (4k)
frame_vm_group_bin_6103 = frame (4k)
frame_vm_group_bin_6104 = frame (4k)
frame_vm_group_bin_6105 = frame (4k)
frame_vm_group_bin_6106 = frame (4k)
frame_vm_group_bin_6107 = frame (4k)
frame_vm_group_bin_6108 = frame (4k)
frame_vm_group_bin_6109 = frame (4k)
frame_vm_group_bin_6110 = frame (4k)
frame_vm_group_bin_6111 = frame (4k)
frame_vm_group_bin_6112 = frame (4k)
frame_vm_group_bin_6113 = frame (4k)
frame_vm_group_bin_6114 = frame (4k)
frame_vm_group_bin_6115 = frame (4k)
frame_vm_group_bin_6116 = frame (4k)
frame_vm_group_bin_6117 = frame (4k)
frame_vm_group_bin_6118 = frame (4k)
frame_vm_group_bin_6119 = frame (4k)
frame_vm_group_bin_6120 = frame (4k)
frame_vm_group_bin_6121 = frame (4k)
frame_vm_group_bin_6122 = frame (4k)
frame_vm_group_bin_6123 = frame (4k)
frame_vm_group_bin_6124 = frame (4k)
frame_vm_group_bin_6125 = frame (4k)
frame_vm_group_bin_6126 = frame (4k)
frame_vm_group_bin_6127 = frame (4k)
frame_vm_group_bin_6128 = frame (4k)
frame_vm_group_bin_6129 = frame (4k)
frame_vm_group_bin_6130 = frame (4k)
frame_vm_group_bin_6131 = frame (4k)
frame_vm_group_bin_6132 = frame (4k)
frame_vm_group_bin_6133 = frame (4k)
frame_vm_group_bin_6134 = frame (4k)
frame_vm_group_bin_6135 = frame (4k)
frame_vm_group_bin_6136 = frame (4k)
frame_vm_group_bin_6137 = frame (4k)
frame_vm_group_bin_6138 = frame (4k)
frame_vm_group_bin_6139 = frame (4k)
frame_vm_group_bin_6140 = frame (4k)
frame_vm_group_bin_6141 = frame (4k)
frame_vm_group_bin_6142 = frame (4k)
frame_vm_group_bin_6143 = frame (4k)
frame_vm_group_bin_6144 = frame (4k)
frame_vm_group_bin_6145 = frame (4k)
frame_vm_group_bin_6146 = frame (4k)
frame_vm_group_bin_6147 = frame (4k)
frame_vm_group_bin_6148 = frame (4k)
frame_vm_group_bin_6149 = frame (4k)
frame_vm_group_bin_6150 = frame (4k)
frame_vm_group_bin_6151 = frame (4k)
frame_vm_group_bin_6152 = frame (4k)
frame_vm_group_bin_6153 = frame (4k)
frame_vm_group_bin_6154 = frame (4k)
frame_vm_group_bin_6155 = frame (4k)
frame_vm_group_bin_6156 = frame (4k)
frame_vm_group_bin_6157 = frame (4k)
frame_vm_group_bin_6158 = frame (4k)
frame_vm_group_bin_6159 = frame (4k)
frame_vm_group_bin_6160 = frame (4k)
frame_vm_group_bin_6161 = frame (4k)
frame_vm_group_bin_6162 = frame (4k)
frame_vm_group_bin_6163 = frame (4k)
frame_vm_group_bin_6164 = frame (4k)
frame_vm_group_bin_6165 = frame (4k)
frame_vm_group_bin_6166 = frame (4k)
frame_vm_group_bin_6167 = frame (4k)
frame_vm_group_bin_6168 = frame (4k)
frame_vm_group_bin_6169 = frame (4k)
frame_vm_group_bin_6170 = frame (4k)
frame_vm_group_bin_6171 = frame (4k)
frame_vm_group_bin_6172 = frame (4k)
frame_vm_group_bin_6173 = frame (4k)
frame_vm_group_bin_6174 = frame (4k)
frame_vm_group_bin_6175 = frame (4k)
frame_vm_group_bin_6176 = frame (4k)
frame_vm_group_bin_6177 = frame (4k)
frame_vm_group_bin_6178 = frame (4k)
frame_vm_group_bin_6179 = frame (4k)
frame_vm_group_bin_6180 = frame (4k)
frame_vm_group_bin_6181 = frame (4k)
frame_vm_group_bin_6182 = frame (4k)
frame_vm_group_bin_6183 = frame (4k)
frame_vm_group_bin_6184 = frame (4k)
frame_vm_group_bin_6185 = frame (4k)
frame_vm_group_bin_6186 = frame (4k)
frame_vm_group_bin_6187 = frame (4k)
frame_vm_group_bin_6188 = frame (4k)
frame_vm_group_bin_6189 = frame (4k)
frame_vm_group_bin_6190 = frame (4k)
frame_vm_group_bin_6191 = frame (4k)
frame_vm_group_bin_6192 = frame (4k)
frame_vm_group_bin_6193 = frame (4k)
frame_vm_group_bin_6194 = frame (4k)
frame_vm_group_bin_6195 = frame (4k)
frame_vm_group_bin_6196 = frame (4k)
frame_vm_group_bin_6197 = frame (4k)
frame_vm_group_bin_6198 = frame (4k)
frame_vm_group_bin_6199 = frame (4k)
frame_vm_group_bin_6200 = frame (4k)
frame_vm_group_bin_6201 = frame (4k)
frame_vm_group_bin_6202 = frame (4k)
frame_vm_group_bin_6203 = frame (4k)
frame_vm_group_bin_6204 = frame (4k)
frame_vm_group_bin_6205 = frame (4k)
frame_vm_group_bin_6206 = frame (4k)
frame_vm_group_bin_6207 = frame (4k)
frame_vm_group_bin_6208 = frame (4k)
frame_vm_group_bin_6209 = frame (4k)
frame_vm_group_bin_6210 = frame (4k)
frame_vm_group_bin_6211 = frame (4k)
frame_vm_group_bin_6212 = frame (4k)
frame_vm_group_bin_6213 = frame (4k)
frame_vm_group_bin_6214 = frame (4k)
frame_vm_group_bin_6215 = frame (4k)
frame_vm_group_bin_6216 = frame (4k)
frame_vm_group_bin_6217 = frame (4k)
frame_vm_group_bin_6218 = frame (4k)
frame_vm_group_bin_6219 = frame (4k)
frame_vm_group_bin_6220 = frame (4k)
frame_vm_group_bin_6221 = frame (4k)
frame_vm_group_bin_6222 = frame (4k)
frame_vm_group_bin_6223 = frame (4k)
frame_vm_group_bin_6224 = frame (4k)
frame_vm_group_bin_6225 = frame (4k)
frame_vm_group_bin_6226 = frame (4k)
frame_vm_group_bin_6227 = frame (4k)
frame_vm_group_bin_6228 = frame (4k)
frame_vm_group_bin_6229 = frame (4k)
frame_vm_group_bin_6230 = frame (4k)
frame_vm_group_bin_6231 = frame (4k)
frame_vm_group_bin_6232 = frame (4k)
frame_vm_group_bin_6233 = frame (4k)
frame_vm_group_bin_6234 = frame (4k)
frame_vm_group_bin_6235 = frame (4k)
frame_vm_group_bin_6236 = frame (4k)
frame_vm_group_bin_6237 = frame (4k)
frame_vm_group_bin_6238 = frame (4k)
frame_vm_group_bin_6239 = frame (4k)
frame_vm_group_bin_6240 = frame (4k)
frame_vm_group_bin_6241 = frame (4k)
frame_vm_group_bin_6242 = frame (4k)
frame_vm_group_bin_6243 = frame (4k)
frame_vm_group_bin_6244 = frame (4k)
frame_vm_group_bin_6245 = frame (4k)
frame_vm_group_bin_6246 = frame (4k)
frame_vm_group_bin_6247 = frame (4k)
frame_vm_group_bin_6248 = frame (4k)
frame_vm_group_bin_6249 = frame (4k)
frame_vm_group_bin_6250 = frame (4k)
frame_vm_group_bin_6251 = frame (4k)
frame_vm_group_bin_6252 = frame (4k)
frame_vm_group_bin_6253 = frame (4k)
frame_vm_group_bin_6254 = frame (4k)
frame_vm_group_bin_6255 = frame (4k)
frame_vm_group_bin_6256 = frame (4k)
frame_vm_group_bin_6257 = frame (4k)
frame_vm_group_bin_6258 = frame (4k)
frame_vm_group_bin_6259 = frame (4k)
frame_vm_group_bin_6260 = frame (4k)
frame_vm_group_bin_6261 = frame (4k)
frame_vm_group_bin_6262 = frame (4k)
frame_vm_group_bin_6263 = frame (4k)
frame_vm_group_bin_6264 = frame (4k)
frame_vm_group_bin_6265 = frame (4k)
frame_vm_group_bin_6266 = frame (4k)
frame_vm_group_bin_6267 = frame (4k)
frame_vm_group_bin_6268 = frame (4k)
frame_vm_group_bin_6269 = frame (4k)
frame_vm_group_bin_6270 = frame (4k)
frame_vm_group_bin_6271 = frame (4k)
frame_vm_group_bin_6272 = frame (4k)
frame_vm_group_bin_6273 = frame (4k)
frame_vm_group_bin_6274 = frame (4k)
frame_vm_group_bin_6275 = frame (4k)
frame_vm_group_bin_6276 = frame (4k)
frame_vm_group_bin_6277 = frame (4k)
frame_vm_group_bin_6278 = frame (4k)
frame_vm_group_bin_6279 = frame (4k)
frame_vm_group_bin_6280 = frame (4k)
frame_vm_group_bin_6281 = frame (4k)
frame_vm_group_bin_6282 = frame (4k)
frame_vm_group_bin_6283 = frame (4k)
frame_vm_group_bin_6284 = frame (4k)
frame_vm_group_bin_6285 = frame (4k)
frame_vm_group_bin_6286 = frame (4k)
frame_vm_group_bin_6287 = frame (4k)
frame_vm_group_bin_6288 = frame (4k)
frame_vm_group_bin_6289 = frame (4k)
frame_vm_group_bin_6290 = frame (4k)
frame_vm_group_bin_6291 = frame (4k)
frame_vm_group_bin_6292 = frame (4k)
frame_vm_group_bin_6293 = frame (4k)
frame_vm_group_bin_6294 = frame (4k)
frame_vm_group_bin_6295 = frame (4k)
frame_vm_group_bin_6296 = frame (4k)
frame_vm_group_bin_6297 = frame (4k)
frame_vm_group_bin_6298 = frame (4k)
frame_vm_group_bin_6299 = frame (4k)
frame_vm_group_bin_6300 = frame (4k)
frame_vm_group_bin_6301 = frame (4k)
frame_vm_group_bin_6302 = frame (4k)
frame_vm_group_bin_6303 = frame (4k)
frame_vm_group_bin_6304 = frame (4k)
frame_vm_group_bin_6305 = frame (4k)
frame_vm_group_bin_6306 = frame (4k)
frame_vm_group_bin_6307 = frame (4k)
frame_vm_group_bin_6308 = frame (4k)
frame_vm_group_bin_6309 = frame (4k)
frame_vm_group_bin_6310 = frame (4k)
frame_vm_group_bin_6311 = frame (4k)
frame_vm_group_bin_6312 = frame (4k)
frame_vm_group_bin_6313 = frame (4k)
frame_vm_group_bin_6314 = frame (4k)
frame_vm_group_bin_6315 = frame (4k)
frame_vm_group_bin_6316 = frame (4k)
frame_vm_group_bin_6317 = frame (4k)
frame_vm_group_bin_6318 = frame (4k)
frame_vm_group_bin_6319 = frame (4k)
frame_vm_group_bin_6320 = frame (4k)
frame_vm_group_bin_6321 = frame (4k)
frame_vm_group_bin_6322 = frame (4k)
frame_vm_group_bin_6323 = frame (4k)
frame_vm_group_bin_6324 = frame (4k)
frame_vm_group_bin_6325 = frame (4k)
frame_vm_group_bin_6326 = frame (4k)
frame_vm_group_bin_6327 = frame (4k)
frame_vm_group_bin_6328 = frame (4k)
frame_vm_group_bin_6329 = frame (4k)
frame_vm_group_bin_6330 = frame (4k)
frame_vm_group_bin_6331 = frame (4k)
frame_vm_group_bin_6332 = frame (4k)
frame_vm_group_bin_6333 = frame (4k)
frame_vm_group_bin_6334 = frame (4k)
frame_vm_group_bin_6335 = frame (4k)
frame_vm_group_bin_6336 = frame (4k)
frame_vm_group_bin_6337 = frame (4k)
frame_vm_group_bin_6338 = frame (4k)
frame_vm_group_bin_6339 = frame (4k)
frame_vm_group_bin_6340 = frame (4k)
frame_vm_group_bin_6341 = frame (4k)
frame_vm_group_bin_6342 = frame (4k)
frame_vm_group_bin_6343 = frame (4k)
frame_vm_group_bin_6344 = frame (4k)
frame_vm_group_bin_6345 = frame (4k)
frame_vm_group_bin_6346 = frame (4k)
frame_vm_group_bin_6347 = frame (4k)
frame_vm_group_bin_6348 = frame (4k)
frame_vm_group_bin_6349 = frame (4k)
frame_vm_group_bin_6350 = frame (4k)
frame_vm_group_bin_6351 = frame (4k)
frame_vm_group_bin_6352 = frame (4k)
frame_vm_group_bin_6353 = frame (4k)
frame_vm_group_bin_6354 = frame (4k)
frame_vm_group_bin_6355 = frame (4k)
frame_vm_group_bin_6356 = frame (4k)
frame_vm_group_bin_6357 = frame (4k)
frame_vm_group_bin_6358 = frame (4k)
frame_vm_group_bin_6359 = frame (4k)
frame_vm_group_bin_6360 = frame (4k)
frame_vm_group_bin_6361 = frame (4k)
frame_vm_group_bin_6362 = frame (4k)
frame_vm_group_bin_6363 = frame (4k)
frame_vm_group_bin_6364 = frame (4k)
frame_vm_group_bin_6365 = frame (4k)
frame_vm_group_bin_6366 = frame (4k)
frame_vm_group_bin_6367 = frame (4k)
frame_vm_group_bin_6368 = frame (4k)
frame_vm_group_bin_6369 = frame (4k)
frame_vm_group_bin_6370 = frame (4k)
frame_vm_group_bin_6371 = frame (4k)
frame_vm_group_bin_6372 = frame (4k)
frame_vm_group_bin_6373 = frame (4k)
frame_vm_group_bin_6374 = frame (4k)
frame_vm_group_bin_6375 = frame (4k)
frame_vm_group_bin_6376 = frame (4k)
frame_vm_group_bin_6377 = frame (4k)
frame_vm_group_bin_6378 = frame (4k)
frame_vm_group_bin_6379 = frame (4k)
frame_vm_group_bin_6380 = frame (4k)
frame_vm_group_bin_6381 = frame (4k)
frame_vm_group_bin_6382 = frame (4k)
frame_vm_group_bin_6383 = frame (4k)
frame_vm_group_bin_6384 = frame (4k)
frame_vm_group_bin_6385 = frame (4k)
frame_vm_group_bin_6386 = frame (4k)
frame_vm_group_bin_6387 = frame (4k)
frame_vm_group_bin_6388 = frame (4k)
frame_vm_group_bin_6389 = frame (4k)
frame_vm_group_bin_6390 = frame (4k)
frame_vm_group_bin_6391 = frame (4k)
frame_vm_group_bin_6392 = frame (4k)
frame_vm_group_bin_6393 = frame (4k)
frame_vm_group_bin_6394 = frame (4k)
frame_vm_group_bin_6395 = frame (4k)
frame_vm_group_bin_6396 = frame (4k)
frame_vm_group_bin_6397 = frame (4k)
frame_vm_group_bin_6398 = frame (4k)
frame_vm_group_bin_6399 = frame (4k)
frame_vm_group_bin_6400 = frame (4k)
frame_vm_group_bin_6401 = frame (4k)
frame_vm_group_bin_6402 = frame (4k)
frame_vm_group_bin_6403 = frame (4k)
frame_vm_group_bin_6404 = frame (4k)
frame_vm_group_bin_6405 = frame (4k)
frame_vm_group_bin_6406 = frame (4k)
frame_vm_group_bin_6407 = frame (4k)
frame_vm_group_bin_6408 = frame (4k)
frame_vm_group_bin_6409 = frame (4k)
frame_vm_group_bin_6410 = frame (4k)
frame_vm_group_bin_6411 = frame (4k)
frame_vm_group_bin_6412 = frame (4k)
frame_vm_group_bin_6413 = frame (4k)
frame_vm_group_bin_6414 = frame (4k)
frame_vm_group_bin_6415 = frame (4k)
frame_vm_group_bin_6416 = frame (4k)
frame_vm_group_bin_6417 = frame (4k)
frame_vm_group_bin_6418 = frame (4k)
frame_vm_group_bin_6419 = frame (4k)
frame_vm_group_bin_6420 = frame (4k)
frame_vm_group_bin_6421 = frame (4k)
frame_vm_group_bin_6422 = frame (4k)
frame_vm_group_bin_6423 = frame (4k)
frame_vm_group_bin_6424 = frame (4k)
frame_vm_group_bin_6425 = frame (4k)
frame_vm_group_bin_6426 = frame (4k)
frame_vm_group_bin_6427 = frame (4k)
frame_vm_group_bin_6428 = frame (4k)
frame_vm_group_bin_6429 = frame (4k)
frame_vm_group_bin_6430 = frame (4k)
frame_vm_group_bin_6431 = frame (4k)
frame_vm_group_bin_6432 = frame (4k)
frame_vm_group_bin_6433 = frame (4k)
frame_vm_group_bin_6434 = frame (4k)
frame_vm_group_bin_6435 = frame (4k)
frame_vm_group_bin_6436 = frame (4k)
frame_vm_group_bin_6437 = frame (4k)
frame_vm_group_bin_6438 = frame (4k)
frame_vm_group_bin_6439 = frame (4k)
frame_vm_group_bin_6440 = frame (4k)
frame_vm_group_bin_6441 = frame (4k)
frame_vm_group_bin_6442 = frame (4k)
frame_vm_group_bin_6443 = frame (4k)
frame_vm_group_bin_6444 = frame (4k)
frame_vm_group_bin_6445 = frame (4k)
frame_vm_group_bin_6446 = frame (4k)
frame_vm_group_bin_6447 = frame (4k)
frame_vm_group_bin_6448 = frame (4k)
frame_vm_group_bin_6449 = frame (4k)
frame_vm_group_bin_6450 = frame (4k)
frame_vm_group_bin_6451 = frame (4k)
frame_vm_group_bin_6452 = frame (4k)
frame_vm_group_bin_6453 = frame (4k)
frame_vm_group_bin_6454 = frame (4k)
frame_vm_group_bin_6455 = frame (4k)
frame_vm_group_bin_6456 = frame (4k)
frame_vm_group_bin_6457 = frame (4k)
frame_vm_group_bin_6458 = frame (4k)
frame_vm_group_bin_6459 = frame (4k)
frame_vm_group_bin_6460 = frame (4k)
frame_vm_group_bin_6461 = frame (4k)
frame_vm_group_bin_6462 = frame (4k)
frame_vm_group_bin_6463 = frame (4k)
frame_vm_group_bin_6464 = frame (4k)
frame_vm_group_bin_6465 = frame (4k)
frame_vm_group_bin_6466 = frame (4k)
frame_vm_group_bin_6467 = frame (4k)
frame_vm_group_bin_6468 = frame (4k)
frame_vm_group_bin_6469 = frame (4k)
frame_vm_group_bin_6470 = frame (4k)
frame_vm_group_bin_6471 = frame (4k)
frame_vm_group_bin_6472 = frame (4k)
frame_vm_group_bin_6473 = frame (4k)
frame_vm_group_bin_6474 = frame (4k)
frame_vm_group_bin_6475 = frame (4k)
frame_vm_group_bin_6476 = frame (4k)
frame_vm_group_bin_6477 = frame (4k)
frame_vm_group_bin_6478 = frame (4k)
frame_vm_group_bin_6479 = frame (4k)
frame_vm_group_bin_6480 = frame (4k)
frame_vm_group_bin_6481 = frame (4k)
frame_vm_group_bin_6482 = frame (4k)
frame_vm_group_bin_6483 = frame (4k)
frame_vm_group_bin_6484 = frame (4k)
frame_vm_group_bin_6485 = frame (4k)
frame_vm_group_bin_6486 = frame (4k)
frame_vm_group_bin_6487 = frame (4k)
frame_vm_group_bin_6488 = frame (4k)
frame_vm_group_bin_6489 = frame (4k)
frame_vm_group_bin_6490 = frame (4k)
frame_vm_group_bin_6491 = frame (4k)
frame_vm_group_bin_6492 = frame (4k)
frame_vm_group_bin_6493 = frame (4k)
frame_vm_group_bin_6494 = frame (4k)
frame_vm_group_bin_6495 = frame (4k)
frame_vm_group_bin_6496 = frame (4k)
frame_vm_group_bin_6497 = frame (4k)
frame_vm_group_bin_6498 = frame (4k)
frame_vm_group_bin_6499 = frame (4k)
frame_vm_group_bin_6500 = frame (4k)
frame_vm_group_bin_6501 = frame (4k)
frame_vm_group_bin_6502 = frame (4k)
frame_vm_group_bin_6503 = frame (4k)
frame_vm_group_bin_6504 = frame (4k)
frame_vm_group_bin_6505 = frame (4k)
frame_vm_group_bin_6506 = frame (4k)
frame_vm_group_bin_6507 = frame (4k)
frame_vm_group_bin_6508 = frame (4k)
frame_vm_group_bin_6509 = frame (4k)
frame_vm_group_bin_6510 = frame (4k)
frame_vm_group_bin_6511 = frame (4k)
frame_vm_group_bin_6512 = frame (4k)
frame_vm_group_bin_6513 = frame (4k)
frame_vm_group_bin_6514 = frame (4k)
frame_vm_group_bin_6515 = frame (4k)
frame_vm_group_bin_6516 = frame (4k)
frame_vm_group_bin_6517 = frame (4k)
frame_vm_group_bin_6518 = frame (4k)
frame_vm_group_bin_6519 = frame (4k)
frame_vm_group_bin_6520 = frame (4k)
frame_vm_group_bin_6521 = frame (4k)
frame_vm_group_bin_6522 = frame (4k)
frame_vm_group_bin_6523 = frame (4k)
frame_vm_group_bin_6524 = frame (4k)
frame_vm_group_bin_6525 = frame (4k)
frame_vm_group_bin_6526 = frame (4k)
frame_vm_group_bin_6527 = frame (4k)
frame_vm_group_bin_6528 = frame (4k)
frame_vm_group_bin_6529 = frame (4k)
frame_vm_group_bin_6530 = frame (4k)
frame_vm_group_bin_6531 = frame (4k)
frame_vm_group_bin_6532 = frame (4k)
frame_vm_group_bin_6533 = frame (4k)
frame_vm_group_bin_6534 = frame (4k)
frame_vm_group_bin_6535 = frame (4k)
frame_vm_group_bin_6536 = frame (4k)
frame_vm_group_bin_6537 = frame (4k)
frame_vm_group_bin_6538 = frame (4k)
frame_vm_group_bin_6539 = frame (4k)
frame_vm_group_bin_6540 = frame (4k)
frame_vm_group_bin_6541 = frame (4k)
frame_vm_group_bin_6542 = frame (4k)
frame_vm_group_bin_6543 = frame (4k)
frame_vm_group_bin_6544 = frame (4k)
frame_vm_group_bin_6545 = frame (4k)
frame_vm_group_bin_6546 = frame (4k)
frame_vm_group_bin_6547 = frame (4k)
frame_vm_group_bin_6548 = frame (4k)
frame_vm_group_bin_6549 = frame (4k)
frame_vm_group_bin_6550 = frame (4k)
frame_vm_group_bin_6551 = frame (4k)
frame_vm_group_bin_6552 = frame (4k)
frame_vm_group_bin_6553 = frame (4k)
frame_vm_group_bin_6554 = frame (4k)
frame_vm_group_bin_6555 = frame (4k)
frame_vm_group_bin_6556 = frame (4k)
frame_vm_group_bin_6557 = frame (4k)
frame_vm_group_bin_6558 = frame (4k)
frame_vm_group_bin_6559 = frame (4k)
frame_vm_group_bin_6560 = frame (4k)
frame_vm_group_bin_6561 = frame (4k)
frame_vm_group_bin_6562 = frame (4k)
frame_vm_group_bin_6563 = frame (4k)
frame_vm_group_bin_6564 = frame (4k)
frame_vm_group_bin_6565 = frame (4k)
frame_vm_group_bin_6566 = frame (4k)
frame_vm_group_bin_6567 = frame (4k)
frame_vm_group_bin_6568 = frame (4k)
frame_vm_group_bin_6569 = frame (4k)
frame_vm_group_bin_6570 = frame (4k)
frame_vm_group_bin_6571 = frame (4k)
frame_vm_group_bin_6572 = frame (4k)
frame_vm_group_bin_6573 = frame (4k)
frame_vm_group_bin_6574 = frame (4k)
frame_vm_group_bin_6575 = frame (4k)
frame_vm_group_bin_6576 = frame (4k)
frame_vm_group_bin_6577 = frame (4k)
frame_vm_group_bin_6578 = frame (4k)
frame_vm_group_bin_6579 = frame (4k)
frame_vm_group_bin_6580 = frame (4k)
frame_vm_group_bin_6581 = frame (4k)
frame_vm_group_bin_6582 = frame (4k)
frame_vm_group_bin_6583 = frame (4k)
frame_vm_group_bin_6584 = frame (4k)
frame_vm_group_bin_6585 = frame (4k)
frame_vm_group_bin_6586 = frame (4k)
frame_vm_group_bin_6587 = frame (4k)
frame_vm_group_bin_6588 = frame (4k)
frame_vm_group_bin_6589 = frame (4k)
frame_vm_group_bin_6590 = frame (4k)
frame_vm_group_bin_6591 = frame (4k)
frame_vm_group_bin_6592 = frame (4k)
frame_vm_group_bin_6593 = frame (4k)
frame_vm_group_bin_6594 = frame (4k)
frame_vm_group_bin_6595 = frame (4k)
frame_vm_group_bin_6596 = frame (4k)
frame_vm_group_bin_6597 = frame (4k)
frame_vm_group_bin_6598 = frame (4k)
frame_vm_group_bin_6599 = frame (4k)
frame_vm_group_bin_6600 = frame (4k)
frame_vm_group_bin_6601 = frame (4k)
frame_vm_group_bin_6602 = frame (4k)
frame_vm_group_bin_6603 = frame (4k)
frame_vm_group_bin_6604 = frame (4k)
frame_vm_group_bin_6605 = frame (4k)
frame_vm_group_bin_6606 = frame (4k)
frame_vm_group_bin_6607 = frame (4k)
frame_vm_group_bin_6608 = frame (4k)
frame_vm_group_bin_6609 = frame (4k)
frame_vm_group_bin_6610 = frame (4k)
frame_vm_group_bin_6611 = frame (4k)
frame_vm_group_bin_6612 = frame (4k)
frame_vm_group_bin_6613 = frame (4k)
frame_vm_group_bin_6614 = frame (4k)
frame_vm_group_bin_6615 = frame (4k)
frame_vm_group_bin_6616 = frame (4k)
frame_vm_group_bin_6617 = frame (4k)
frame_vm_group_bin_6618 = frame (4k)
frame_vm_group_bin_6619 = frame (4k)
frame_vm_group_bin_6620 = frame (4k)
frame_vm_group_bin_6621 = frame (4k)
frame_vm_group_bin_6622 = frame (4k)
frame_vm_group_bin_6623 = frame (4k)
frame_vm_group_bin_6624 = frame (4k)
frame_vm_group_bin_6625 = frame (4k)
frame_vm_group_bin_6626 = frame (4k)
frame_vm_group_bin_6627 = frame (4k)
frame_vm_group_bin_6628 = frame (4k)
frame_vm_group_bin_6629 = frame (4k)
frame_vm_group_bin_6630 = frame (4k)
frame_vm_group_bin_6631 = frame (4k)
frame_vm_group_bin_6632 = frame (4k)
frame_vm_group_bin_6633 = frame (4k)
frame_vm_group_bin_6634 = frame (4k)
frame_vm_group_bin_6635 = frame (4k)
frame_vm_group_bin_6636 = frame (4k)
frame_vm_group_bin_6637 = frame (4k)
frame_vm_group_bin_6638 = frame (4k)
frame_vm_group_bin_6639 = frame (4k)
frame_vm_group_bin_6640 = frame (4k)
frame_vm_group_bin_6641 = frame (4k)
frame_vm_group_bin_6642 = frame (4k)
frame_vm_group_bin_6643 = frame (4k)
frame_vm_group_bin_6644 = frame (4k)
frame_vm_group_bin_6645 = frame (4k)
frame_vm_group_bin_6646 = frame (4k)
frame_vm_group_bin_6647 = frame (4k)
frame_vm_group_bin_6648 = frame (4k)
frame_vm_group_bin_6649 = frame (4k)
frame_vm_group_bin_6650 = frame (4k)
frame_vm_group_bin_6651 = frame (4k)
frame_vm_group_bin_6652 = frame (4k)
frame_vm_group_bin_6653 = frame (4k)
frame_vm_group_bin_6654 = frame (4k)
frame_vm_group_bin_6655 = frame (4k)
frame_vm_group_bin_6656 = frame (4k)
frame_vm_group_bin_6657 = frame (4k)
frame_vm_group_bin_6658 = frame (4k)
frame_vm_group_bin_6659 = frame (4k)
frame_vm_group_bin_6660 = frame (4k)
frame_vm_group_bin_6661 = frame (4k)
frame_vm_group_bin_6662 = frame (4k)
frame_vm_group_bin_6663 = frame (4k)
frame_vm_group_bin_6664 = frame (4k)
frame_vm_group_bin_6665 = frame (4k)
frame_vm_group_bin_6666 = frame (4k)
frame_vm_group_bin_6667 = frame (4k)
frame_vm_group_bin_6668 = frame (4k)
frame_vm_group_bin_6669 = frame (4k)
frame_vm_group_bin_6670 = frame (4k)
frame_vm_group_bin_6671 = frame (4k)
frame_vm_group_bin_6672 = frame (4k)
frame_vm_group_bin_6673 = frame (4k)
frame_vm_group_bin_6674 = frame (4k)
frame_vm_group_bin_6675 = frame (4k)
frame_vm_group_bin_6676 = frame (4k)
frame_vm_group_bin_6677 = frame (4k)
frame_vm_group_bin_6678 = frame (4k)
frame_vm_group_bin_6679 = frame (4k)
frame_vm_group_bin_6680 = frame (4k)
frame_vm_group_bin_6681 = frame (4k)
frame_vm_group_bin_6682 = frame (4k)
frame_vm_group_bin_6683 = frame (4k)
frame_vm_group_bin_6684 = frame (4k)
frame_vm_group_bin_6685 = frame (4k)
frame_vm_group_bin_6686 = frame (4k)
frame_vm_group_bin_6687 = frame (4k)
frame_vm_group_bin_6688 = frame (4k)
frame_vm_group_bin_6689 = frame (4k)
frame_vm_group_bin_6690 = frame (4k)
frame_vm_group_bin_6691 = frame (4k)
frame_vm_group_bin_6692 = frame (4k)
frame_vm_group_bin_6693 = frame (4k)
frame_vm_group_bin_6694 = frame (4k)
frame_vm_group_bin_6695 = frame (4k)
frame_vm_group_bin_6696 = frame (4k)
frame_vm_group_bin_6697 = frame (4k)
frame_vm_group_bin_6698 = frame (4k)
frame_vm_group_bin_6699 = frame (4k)
frame_vm_group_bin_6700 = frame (4k)
frame_vm_group_bin_6701 = frame (4k)
frame_vm_group_bin_6702 = frame (4k)
frame_vm_group_bin_6703 = frame (4k)
frame_vm_group_bin_6704 = frame (4k)
frame_vm_group_bin_6705 = frame (4k)
frame_vm_group_bin_6706 = frame (4k)
frame_vm_group_bin_6707 = frame (4k)
frame_vm_group_bin_6708 = frame (4k)
frame_vm_group_bin_6709 = frame (4k)
frame_vm_group_bin_6710 = frame (4k)
frame_vm_group_bin_6711 = frame (4k)
frame_vm_group_bin_6712 = frame (4k)
frame_vm_group_bin_6713 = frame (4k)
frame_vm_group_bin_6714 = frame (4k)
frame_vm_group_bin_6715 = frame (4k)
frame_vm_group_bin_6716 = frame (4k)
frame_vm_group_bin_6717 = frame (4k)
frame_vm_group_bin_6718 = frame (4k)
frame_vm_group_bin_6719 = frame (4k)
frame_vm_group_bin_6720 = frame (4k)
frame_vm_group_bin_6721 = frame (4k)
frame_vm_group_bin_6722 = frame (4k)
frame_vm_group_bin_6723 = frame (4k)
frame_vm_group_bin_6724 = frame (4k)
frame_vm_group_bin_6725 = frame (4k)
frame_vm_group_bin_6726 = frame (4k)
frame_vm_group_bin_6727 = frame (4k)
frame_vm_group_bin_6728 = frame (4k)
frame_vm_group_bin_6729 = frame (4k)
frame_vm_group_bin_6730 = frame (4k)
frame_vm_group_bin_6731 = frame (4k)
frame_vm_group_bin_6732 = frame (4k)
frame_vm_group_bin_6733 = frame (4k)
frame_vm_group_bin_6734 = frame (4k)
frame_vm_group_bin_6735 = frame (4k)
frame_vm_group_bin_6736 = frame (4k)
frame_vm_group_bin_6737 = frame (4k)
frame_vm_group_bin_6738 = frame (4k)
frame_vm_group_bin_6739 = frame (4k)
frame_vm_group_bin_6740 = frame (4k)
frame_vm_group_bin_6741 = frame (4k)
frame_vm_group_bin_6742 = frame (4k)
frame_vm_group_bin_6743 = frame (4k)
frame_vm_group_bin_6744 = frame (4k)
frame_vm_group_bin_6745 = frame (4k)
frame_vm_group_bin_6746 = frame (4k)
frame_vm_group_bin_6747 = frame (4k)
frame_vm_group_bin_6748 = frame (4k)
frame_vm_group_bin_6749 = frame (4k)
frame_vm_group_bin_6750 = frame (4k)
frame_vm_group_bin_6751 = frame (4k)
frame_vm_group_bin_6752 = frame (4k)
frame_vm_group_bin_6753 = frame (4k)
frame_vm_group_bin_6754 = frame (4k)
frame_vm_group_bin_6755 = frame (4k)
frame_vm_group_bin_6756 = frame (4k)
frame_vm_group_bin_6757 = frame (4k)
frame_vm_group_bin_6758 = frame (4k)
frame_vm_group_bin_6759 = frame (4k)
frame_vm_group_bin_6760 = frame (4k)
frame_vm_group_bin_6761 = frame (4k)
frame_vm_group_bin_6762 = frame (4k)
frame_vm_group_bin_6763 = frame (4k)
frame_vm_group_bin_6764 = frame (4k)
frame_vm_group_bin_6765 = frame (4k)
frame_vm_group_bin_6766 = frame (4k)
frame_vm_group_bin_6767 = frame (4k)
frame_vm_group_bin_6768 = frame (4k)
frame_vm_group_bin_6769 = frame (4k)
frame_vm_group_bin_6770 = frame (4k)
frame_vm_group_bin_6771 = frame (4k)
frame_vm_group_bin_6772 = frame (4k)
frame_vm_group_bin_6773 = frame (4k)
frame_vm_group_bin_6774 = frame (4k)
frame_vm_group_bin_6775 = frame (4k)
frame_vm_group_bin_6776 = frame (4k)
frame_vm_group_bin_6777 = frame (4k)
frame_vm_group_bin_6778 = frame (4k)
frame_vm_group_bin_6779 = frame (4k)
frame_vm_group_bin_6780 = frame (4k)
frame_vm_group_bin_6781 = frame (4k)
frame_vm_group_bin_6782 = frame (4k)
frame_vm_group_bin_6783 = frame (4k)
frame_vm_group_bin_6784 = frame (4k)
frame_vm_group_bin_6785 = frame (4k)
frame_vm_group_bin_6786 = frame (4k)
frame_vm_group_bin_6787 = frame (4k)
frame_vm_group_bin_6788 = frame (4k)
frame_vm_group_bin_6789 = frame (4k)
frame_vm_group_bin_6790 = frame (4k)
frame_vm_group_bin_6791 = frame (4k)
frame_vm_group_bin_6792 = frame (4k)
frame_vm_group_bin_6793 = frame (4k)
frame_vm_group_bin_6794 = frame (4k)
frame_vm_group_bin_6795 = frame (4k)
frame_vm_group_bin_6796 = frame (4k)
frame_vm_group_bin_6797 = frame (4k)
frame_vm_group_bin_6798 = frame (4k)
frame_vm_group_bin_6799 = frame (4k)
frame_vm_group_bin_6800 = frame (4k)
frame_vm_group_bin_6801 = frame (4k)
frame_vm_group_bin_6802 = frame (4k)
frame_vm_group_bin_6803 = frame (4k)
frame_vm_group_bin_6804 = frame (4k)
frame_vm_group_bin_6805 = frame (4k)
frame_vm_group_bin_6806 = frame (4k)
frame_vm_group_bin_6807 = frame (4k)
frame_vm_group_bin_6808 = frame (4k)
frame_vm_group_bin_6809 = frame (4k)
frame_vm_group_bin_6810 = frame (4k)
frame_vm_group_bin_6811 = frame (4k)
frame_vm_group_bin_6812 = frame (4k)
frame_vm_group_bin_6813 = frame (4k)
frame_vm_group_bin_6814 = frame (4k)
frame_vm_group_bin_6815 = frame (4k)
frame_vm_group_bin_6816 = frame (4k)
frame_vm_group_bin_6817 = frame (4k)
frame_vm_group_bin_6818 = frame (4k)
frame_vm_group_bin_6819 = frame (4k)
frame_vm_group_bin_6820 = frame (4k)
frame_vm_group_bin_6821 = frame (4k)
frame_vm_group_bin_6822 = frame (4k)
frame_vm_group_bin_6823 = frame (4k)
frame_vm_group_bin_6824 = frame (4k)
frame_vm_group_bin_6825 = frame (4k)
frame_vm_group_bin_6826 = frame (4k)
frame_vm_group_bin_6827 = frame (4k)
frame_vm_group_bin_6828 = frame (4k)
frame_vm_group_bin_6829 = frame (4k)
frame_vm_group_bin_6830 = frame (4k)
frame_vm_group_bin_6831 = frame (4k)
frame_vm_group_bin_6832 = frame (4k)
frame_vm_group_bin_6833 = frame (4k)
frame_vm_group_bin_6834 = frame (4k)
frame_vm_group_bin_6835 = frame (4k)
frame_vm_group_bin_6836 = frame (4k)
frame_vm_group_bin_6837 = frame (4k)
frame_vm_group_bin_6838 = frame (4k)
frame_vm_group_bin_6839 = frame (4k)
frame_vm_group_bin_6840 = frame (4k)
frame_vm_group_bin_6841 = frame (4k)
frame_vm_group_bin_6842 = frame (4k)
frame_vm_group_bin_6843 = frame (4k)
frame_vm_group_bin_6844 = frame (4k)
frame_vm_group_bin_6845 = frame (4k)
frame_vm_group_bin_6846 = frame (4k)
frame_vm_group_bin_6847 = frame (4k)
frame_vm_group_bin_6848 = frame (4k)
frame_vm_group_bin_6849 = frame (4k)
frame_vm_group_bin_6850 = frame (4k)
frame_vm_group_bin_6851 = frame (4k)
frame_vm_group_bin_6852 = frame (4k)
frame_vm_group_bin_6853 = frame (4k)
frame_vm_group_bin_6854 = frame (4k)
frame_vm_group_bin_6855 = frame (4k)
frame_vm_group_bin_6856 = frame (4k)
frame_vm_group_bin_6857 = frame (4k)
frame_vm_group_bin_6858 = frame (4k)
frame_vm_group_bin_6859 = frame (4k)
frame_vm_group_bin_6860 = frame (4k)
frame_vm_group_bin_6861 = frame (4k)
frame_vm_group_bin_6862 = frame (4k)
frame_vm_group_bin_6863 = frame (4k)
frame_vm_group_bin_6864 = frame (4k)
frame_vm_group_bin_6865 = frame (4k)
frame_vm_group_bin_6866 = frame (4k)
frame_vm_group_bin_6867 = frame (4k)
frame_vm_group_bin_6868 = frame (4k)
frame_vm_group_bin_6869 = frame (4k)
frame_vm_group_bin_6870 = frame (4k)
frame_vm_group_bin_6871 = frame (4k)
frame_vm_group_bin_6872 = frame (4k)
frame_vm_group_bin_6873 = frame (4k)
frame_vm_group_bin_6874 = frame (4k)
frame_vm_group_bin_6875 = frame (4k)
frame_vm_group_bin_6876 = frame (4k)
frame_vm_group_bin_6877 = frame (4k)
frame_vm_group_bin_6878 = frame (4k)
frame_vm_group_bin_6879 = frame (4k)
frame_vm_group_bin_6880 = frame (4k)
frame_vm_group_bin_6881 = frame (4k)
frame_vm_group_bin_6882 = frame (4k)
frame_vm_group_bin_6883 = frame (4k)
frame_vm_group_bin_6884 = frame (4k)
frame_vm_group_bin_6885 = frame (4k)
frame_vm_group_bin_6886 = frame (4k)
frame_vm_group_bin_6887 = frame (4k)
frame_vm_group_bin_6888 = frame (4k)
frame_vm_group_bin_6889 = frame (4k)
frame_vm_group_bin_6890 = frame (4k)
frame_vm_group_bin_6891 = frame (4k)
frame_vm_group_bin_6892 = frame (4k)
frame_vm_group_bin_6893 = frame (4k)
frame_vm_group_bin_6894 = frame (4k)
frame_vm_group_bin_6895 = frame (4k)
frame_vm_group_bin_6896 = frame (4k)
frame_vm_group_bin_6897 = frame (4k)
frame_vm_group_bin_6898 = frame (4k)
frame_vm_group_bin_6899 = frame (4k)
frame_vm_group_bin_6900 = frame (4k)
frame_vm_group_bin_6901 = frame (4k)
frame_vm_group_bin_6902 = frame (4k)
frame_vm_group_bin_6903 = frame (4k)
frame_vm_group_bin_6904 = frame (4k)
frame_vm_group_bin_6905 = frame (4k)
frame_vm_group_bin_6906 = frame (4k)
frame_vm_group_bin_6907 = frame (4k)
frame_vm_group_bin_6908 = frame (4k)
frame_vm_group_bin_6909 = frame (4k)
frame_vm_group_bin_6910 = frame (4k)
frame_vm_group_bin_6911 = frame (4k)
frame_vm_group_bin_6912 = frame (4k)
frame_vm_group_bin_6913 = frame (4k)
frame_vm_group_bin_6914 = frame (4k)
frame_vm_group_bin_6915 = frame (4k)
frame_vm_group_bin_6916 = frame (4k)
frame_vm_group_bin_6917 = frame (4k)
frame_vm_group_bin_6918 = frame (4k)
frame_vm_group_bin_6919 = frame (4k)
frame_vm_group_bin_6920 = frame (4k)
frame_vm_group_bin_6921 = frame (4k)
frame_vm_group_bin_6922 = frame (4k)
frame_vm_group_bin_6923 = frame (4k)
frame_vm_group_bin_6924 = frame (4k)
frame_vm_group_bin_6925 = frame (4k)
frame_vm_group_bin_6926 = frame (4k)
frame_vm_group_bin_6927 = frame (4k)
frame_vm_group_bin_6928 = frame (4k)
frame_vm_group_bin_6929 = frame (4k)
frame_vm_group_bin_6930 = frame (4k)
frame_vm_group_bin_6931 = frame (4k)
frame_vm_group_bin_6932 = frame (4k)
frame_vm_group_bin_6933 = frame (4k)
frame_vm_group_bin_6934 = frame (4k)
frame_vm_group_bin_6935 = frame (4k)
frame_vm_group_bin_6936 = frame (4k)
frame_vm_group_bin_6937 = frame (4k)
frame_vm_group_bin_6938 = frame (4k)
frame_vm_group_bin_6939 = frame (4k)
frame_vm_group_bin_6940 = frame (4k)
frame_vm_group_bin_6941 = frame (4k)
frame_vm_group_bin_6942 = frame (4k)
frame_vm_group_bin_6943 = frame (4k)
frame_vm_group_bin_6944 = frame (4k)
frame_vm_group_bin_6945 = frame (4k)
frame_vm_group_bin_6946 = frame (4k)
frame_vm_group_bin_6947 = frame (4k)
frame_vm_group_bin_6948 = frame (4k)
frame_vm_group_bin_6949 = frame (4k)
frame_vm_group_bin_6950 = frame (4k)
frame_vm_group_bin_6951 = frame (4k)
frame_vm_group_bin_6952 = frame (4k)
frame_vm_group_bin_6953 = frame (4k)
frame_vm_group_bin_6954 = frame (4k)
frame_vm_group_bin_6955 = frame (4k)
frame_vm_group_bin_6956 = frame (4k)
frame_vm_group_bin_6957 = frame (4k)
frame_vm_group_bin_6958 = frame (4k)
frame_vm_group_bin_6959 = frame (4k)
frame_vm_group_bin_6960 = frame (4k)
frame_vm_group_bin_6961 = frame (4k)
frame_vm_group_bin_6962 = frame (4k)
frame_vm_group_bin_6963 = frame (4k)
frame_vm_group_bin_6964 = frame (4k)
frame_vm_group_bin_6965 = frame (4k)
frame_vm_group_bin_6966 = frame (4k)
frame_vm_group_bin_6967 = frame (4k)
frame_vm_group_bin_6968 = frame (4k)
frame_vm_group_bin_6969 = frame (4k)
frame_vm_group_bin_6970 = frame (4k)
frame_vm_group_bin_6971 = frame (4k)
frame_vm_group_bin_6972 = frame (4k)
frame_vm_group_bin_6973 = frame (4k)
frame_vm_group_bin_6974 = frame (4k)
frame_vm_group_bin_6975 = frame (4k)
frame_vm_group_bin_6976 = frame (4k)
frame_vm_group_bin_6977 = frame (4k)
frame_vm_group_bin_6978 = frame (4k)
frame_vm_group_bin_6979 = frame (4k)
frame_vm_group_bin_6980 = frame (4k)
frame_vm_group_bin_6981 = frame (4k)
frame_vm_group_bin_6982 = frame (4k)
frame_vm_group_bin_6983 = frame (4k)
frame_vm_group_bin_6984 = frame (4k)
frame_vm_group_bin_6985 = frame (4k)
frame_vm_group_bin_6986 = frame (4k)
frame_vm_group_bin_6987 = frame (4k)
frame_vm_group_bin_6988 = frame (4k)
frame_vm_group_bin_6989 = frame (4k)
frame_vm_group_bin_6990 = frame (4k)
frame_vm_group_bin_6991 = frame (4k)
frame_vm_group_bin_6992 = frame (4k)
frame_vm_group_bin_6993 = frame (4k)
frame_vm_group_bin_6994 = frame (4k)
frame_vm_group_bin_6995 = frame (4k)
frame_vm_group_bin_6996 = frame (4k)
frame_vm_group_bin_6997 = frame (4k)
frame_vm_group_bin_6998 = frame (4k)
frame_vm_group_bin_6999 = frame (4k)
frame_vm_group_bin_7000 = frame (4k)
frame_vm_group_bin_7001 = frame (4k)
frame_vm_group_bin_7002 = frame (4k)
frame_vm_group_bin_7003 = frame (4k)
frame_vm_group_bin_7004 = frame (4k)
frame_vm_group_bin_7005 = frame (4k)
frame_vm_group_bin_7006 = frame (4k)
frame_vm_group_bin_7007 = frame (4k)
frame_vm_group_bin_7008 = frame (4k)
frame_vm_group_bin_7009 = frame (4k)
frame_vm_group_bin_7010 = frame (4k)
frame_vm_group_bin_7011 = frame (4k)
frame_vm_group_bin_7012 = frame (4k)
frame_vm_group_bin_7013 = frame (4k)
frame_vm_group_bin_7014 = frame (4k)
frame_vm_group_bin_7015 = frame (4k)
frame_vm_group_bin_7016 = frame (4k)
frame_vm_group_bin_7017 = frame (4k)
frame_vm_group_bin_7018 = frame (4k)
frame_vm_group_bin_7019 = frame (4k)
frame_vm_group_bin_7020 = frame (4k)
frame_vm_group_bin_7021 = frame (4k)
frame_vm_group_bin_7022 = frame (4k)
frame_vm_group_bin_7023 = frame (4k)
frame_vm_group_bin_7024 = frame (4k)
frame_vm_group_bin_7025 = frame (4k)
frame_vm_group_bin_7026 = frame (4k)
frame_vm_group_bin_7027 = frame (4k)
frame_vm_group_bin_7028 = frame (4k)
frame_vm_group_bin_7029 = frame (4k)
frame_vm_group_bin_7030 = frame (4k)
frame_vm_group_bin_7031 = frame (4k)
frame_vm_group_bin_7032 = frame (4k)
frame_vm_group_bin_7033 = frame (4k)
frame_vm_group_bin_7034 = frame (4k)
frame_vm_group_bin_7035 = frame (4k)
frame_vm_group_bin_7036 = frame (4k)
frame_vm_group_bin_7037 = frame (4k)
frame_vm_group_bin_7038 = frame (4k)
frame_vm_group_bin_7039 = frame (4k)
frame_vm_group_bin_7040 = frame (4k)
frame_vm_group_bin_7041 = frame (4k)
frame_vm_group_bin_7042 = frame (4k)
frame_vm_group_bin_7043 = frame (4k)
frame_vm_group_bin_7044 = frame (4k)
frame_vm_group_bin_7045 = frame (4k)
frame_vm_group_bin_7046 = frame (4k)
frame_vm_group_bin_7047 = frame (4k)
frame_vm_group_bin_7048 = frame (4k)
frame_vm_group_bin_7049 = frame (4k)
frame_vm_group_bin_7050 = frame (4k)
frame_vm_group_bin_7051 = frame (4k)
frame_vm_group_bin_7052 = frame (4k)
frame_vm_group_bin_7053 = frame (4k)
frame_vm_group_bin_7054 = frame (4k)
frame_vm_group_bin_7055 = frame (4k)
frame_vm_group_bin_7056 = frame (4k)
frame_vm_group_bin_7057 = frame (4k)
frame_vm_group_bin_7058 = frame (4k)
frame_vm_group_bin_7059 = frame (4k)
frame_vm_group_bin_7060 = frame (4k)
frame_vm_group_bin_7061 = frame (4k)
frame_vm_group_bin_7062 = frame (4k)
frame_vm_group_bin_7063 = frame (4k)
frame_vm_group_bin_7064 = frame (4k)
frame_vm_group_bin_7065 = frame (4k)
frame_vm_group_bin_7066 = frame (4k)
frame_vm_group_bin_7067 = frame (4k)
frame_vm_group_bin_7068 = frame (4k)
frame_vm_group_bin_7069 = frame (4k)
frame_vm_group_bin_7070 = frame (4k)
frame_vm_group_bin_7071 = frame (4k)
frame_vm_group_bin_7072 = frame (4k)
frame_vm_group_bin_7073 = frame (4k)
frame_vm_group_bin_7074 = frame (4k)
frame_vm_group_bin_7075 = frame (4k)
frame_vm_group_bin_7076 = frame (4k)
frame_vm_group_bin_7077 = frame (4k)
frame_vm_group_bin_7078 = frame (4k)
frame_vm_group_bin_7079 = frame (4k)
frame_vm_group_bin_7080 = frame (4k)
frame_vm_group_bin_7081 = frame (4k)
frame_vm_group_bin_7082 = frame (4k)
frame_vm_group_bin_7083 = frame (4k)
frame_vm_group_bin_7084 = frame (4k)
frame_vm_group_bin_7085 = frame (4k)
frame_vm_group_bin_7086 = frame (4k)
frame_vm_group_bin_7087 = frame (4k)
frame_vm_group_bin_7088 = frame (4k)
frame_vm_group_bin_7089 = frame (4k)
frame_vm_group_bin_7090 = frame (4k)
frame_vm_group_bin_7091 = frame (4k)
frame_vm_group_bin_7092 = frame (4k)
frame_vm_group_bin_7093 = frame (4k)
frame_vm_group_bin_7094 = frame (4k)
frame_vm_group_bin_7095 = frame (4k)
frame_vm_group_bin_7096 = frame (4k)
frame_vm_group_bin_7097 = frame (4k)
frame_vm_group_bin_7098 = frame (4k)
frame_vm_group_bin_7099 = frame (4k)
frame_vm_group_bin_7100 = frame (4k)
frame_vm_group_bin_7101 = frame (4k)
frame_vm_group_bin_7102 = frame (4k)
frame_vm_group_bin_7103 = frame (4k)
frame_vm_group_bin_7104 = frame (4k)
frame_vm_group_bin_7105 = frame (4k)
frame_vm_group_bin_7106 = frame (4k)
frame_vm_group_bin_7107 = frame (4k)
frame_vm_group_bin_7108 = frame (4k)
frame_vm_group_bin_7109 = frame (4k)
frame_vm_group_bin_7110 = frame (4k)
frame_vm_group_bin_7111 = frame (4k)
frame_vm_group_bin_7112 = frame (4k)
frame_vm_group_bin_7113 = frame (4k)
frame_vm_group_bin_7114 = frame (4k)
frame_vm_group_bin_7115 = frame (4k)
frame_vm_group_bin_7116 = frame (4k)
frame_vm_group_bin_7117 = frame (4k)
frame_vm_group_bin_7118 = frame (4k)
frame_vm_group_bin_7119 = frame (4k)
frame_vm_group_bin_7120 = frame (4k)
frame_vm_group_bin_7121 = frame (4k)
frame_vm_group_bin_7122 = frame (4k)
frame_vm_group_bin_7123 = frame (4k)
frame_vm_group_bin_7124 = frame (4k)
frame_vm_group_bin_7125 = frame (4k)
frame_vm_group_bin_7126 = frame (4k)
frame_vm_group_bin_7127 = frame (4k)
frame_vm_group_bin_7128 = frame (4k)
frame_vm_group_bin_7129 = frame (4k)
frame_vm_group_bin_7130 = frame (4k)
frame_vm_group_bin_7131 = frame (4k)
frame_vm_group_bin_7132 = frame (4k)
frame_vm_group_bin_7133 = frame (4k)
frame_vm_group_bin_7134 = frame (4k)
frame_vm_group_bin_7135 = frame (4k)
frame_vm_group_bin_7136 = frame (4k)
frame_vm_group_bin_7137 = frame (4k)
frame_vm_group_bin_7138 = frame (4k)
frame_vm_group_bin_7139 = frame (4k)
frame_vm_group_bin_7140 = frame (4k)
frame_vm_group_bin_7141 = frame (4k)
frame_vm_group_bin_7142 = frame (4k)
frame_vm_group_bin_7143 = frame (4k)
frame_vm_group_bin_7144 = frame (4k)
frame_vm_group_bin_7145 = frame (4k)
frame_vm_group_bin_7146 = frame (4k)
frame_vm_group_bin_7147 = frame (4k)
frame_vm_group_bin_7148 = frame (4k)
frame_vm_group_bin_7149 = frame (4k)
frame_vm_group_bin_7150 = frame (4k)
frame_vm_group_bin_7151 = frame (4k)
frame_vm_group_bin_7152 = frame (4k)
frame_vm_group_bin_7153 = frame (4k)
frame_vm_group_bin_7154 = frame (4k)
frame_vm_group_bin_7155 = frame (4k)
frame_vm_group_bin_7156 = frame (4k)
frame_vm_group_bin_7157 = frame (4k)
frame_vm_group_bin_7158 = frame (4k)
frame_vm_group_bin_7159 = frame (4k)
frame_vm_group_bin_7160 = frame (4k)
frame_vm_group_bin_7161 = frame (4k)
frame_vm_group_bin_7162 = frame (4k)
frame_vm_group_bin_7163 = frame (4k)
frame_vm_group_bin_7164 = frame (4k)
frame_vm_group_bin_7165 = frame (4k)
frame_vm_group_bin_7166 = frame (4k)
frame_vm_group_bin_7167 = frame (4k)
frame_vm_group_bin_7168 = frame (4k)
frame_vm_group_bin_7169 = frame (4k)
frame_vm_group_bin_7170 = frame (4k)
frame_vm_group_bin_7171 = frame (4k)
frame_vm_group_bin_7172 = frame (4k)
frame_vm_group_bin_7173 = frame (4k)
frame_vm_group_bin_7174 = frame (4k)
frame_vm_group_bin_7175 = frame (4k)
frame_vm_group_bin_7176 = frame (4k)
frame_vm_group_bin_7177 = frame (4k)
frame_vm_group_bin_7178 = frame (4k)
frame_vm_group_bin_7179 = frame (4k)
frame_vm_group_bin_7180 = frame (4k)
frame_vm_group_bin_7181 = frame (4k)
frame_vm_group_bin_7182 = frame (4k)
frame_vm_group_bin_7183 = frame (4k)
frame_vm_group_bin_7184 = frame (4k)
frame_vm_group_bin_7185 = frame (4k)
frame_vm_group_bin_7186 = frame (4k)
frame_vm_group_bin_7187 = frame (4k)
frame_vm_group_bin_7188 = frame (4k)
frame_vm_group_bin_7189 = frame (4k)
frame_vm_group_bin_7190 = frame (4k)
frame_vm_group_bin_7191 = frame (4k)
frame_vm_group_bin_7192 = frame (4k)
frame_vm_group_bin_7193 = frame (4k)
frame_vm_group_bin_7194 = frame (4k)
frame_vm_group_bin_7195 = frame (4k)
frame_vm_group_bin_7196 = frame (4k)
frame_vm_group_bin_7197 = frame (4k)
frame_vm_group_bin_7198 = frame (4k)
frame_vm_group_bin_7199 = frame (4k)
frame_vm_group_bin_7200 = frame (4k)
frame_vm_group_bin_7201 = frame (4k)
frame_vm_group_bin_7202 = frame (4k)
frame_vm_group_bin_7203 = frame (4k)
frame_vm_group_bin_7204 = frame (4k)
frame_vm_group_bin_7205 = frame (4k)
frame_vm_group_bin_7206 = frame (4k)
frame_vm_group_bin_7207 = frame (4k)
frame_vm_group_bin_7208 = frame (4k)
frame_vm_group_bin_7209 = frame (4k)
frame_vm_group_bin_7210 = frame (4k)
frame_vm_group_bin_7211 = frame (4k)
frame_vm_group_bin_7212 = frame (4k)
frame_vm_group_bin_7213 = frame (4k)
frame_vm_group_bin_7214 = frame (4k)
frame_vm_group_bin_7215 = frame (4k)
frame_vm_group_bin_7216 = frame (4k)
frame_vm_group_bin_7217 = frame (4k)
frame_vm_group_bin_7218 = frame (4k)
frame_vm_group_bin_7219 = frame (4k)
frame_vm_group_bin_7220 = frame (4k)
frame_vm_group_bin_7221 = frame (4k)
frame_vm_group_bin_7222 = frame (4k)
frame_vm_group_bin_7223 = frame (4k)
frame_vm_group_bin_7224 = frame (4k)
frame_vm_group_bin_7225 = frame (4k)
frame_vm_group_bin_7226 = frame (4k)
frame_vm_group_bin_7227 = frame (4k)
frame_vm_group_bin_7228 = frame (4k)
frame_vm_group_bin_7229 = frame (4k)
frame_vm_group_bin_7230 = frame (4k)
frame_vm_group_bin_7231 = frame (4k)
frame_vm_group_bin_7232 = frame (4k)
frame_vm_group_bin_7233 = frame (4k)
frame_vm_group_bin_7234 = frame (4k)
frame_vm_group_bin_7235 = frame (4k)
frame_vm_group_bin_7236 = frame (4k)
frame_vm_group_bin_7237 = frame (4k)
frame_vm_group_bin_7238 = frame (4k)
frame_vm_group_bin_7239 = frame (4k)
frame_vm_group_bin_7240 = frame (4k)
frame_vm_group_bin_7241 = frame (4k)
frame_vm_group_bin_7242 = frame (4k)
frame_vm_group_bin_7243 = frame (4k)
frame_vm_group_bin_7244 = frame (4k)
frame_vm_group_bin_7245 = frame (4k)
frame_vm_group_bin_7246 = frame (4k)
frame_vm_group_bin_7247 = frame (4k)
frame_vm_group_bin_7248 = frame (4k)
frame_vm_group_bin_7249 = frame (4k)
frame_vm_group_bin_7250 = frame (4k)
frame_vm_group_bin_7251 = frame (4k)
frame_vm_group_bin_7252 = frame (4k)
frame_vm_group_bin_7253 = frame (4k)
frame_vm_group_bin_7254 = frame (4k)
frame_vm_group_bin_7255 = frame (4k)
frame_vm_group_bin_7256 = frame (4k)
frame_vm_group_bin_7257 = frame (4k)
frame_vm_group_bin_7258 = frame (4k)
frame_vm_group_bin_7259 = frame (4k)
frame_vm_group_bin_7260 = frame (4k)
frame_vm_group_bin_7261 = frame (4k)
frame_vm_group_bin_7262 = frame (4k)
frame_vm_group_bin_7263 = frame (4k)
frame_vm_group_bin_7264 = frame (4k)
frame_vm_group_bin_7265 = frame (4k)
frame_vm_group_bin_7266 = frame (4k)
frame_vm_group_bin_7267 = frame (4k)
frame_vm_group_bin_7268 = frame (4k)
frame_vm_group_bin_7269 = frame (4k)
frame_vm_group_bin_7270 = frame (4k)
frame_vm_group_bin_7271 = frame (4k)
frame_vm_group_bin_7272 = frame (4k)
frame_vm_group_bin_7273 = frame (4k)
frame_vm_group_bin_7274 = frame (4k)
frame_vm_group_bin_7275 = frame (4k)
frame_vm_group_bin_7276 = frame (4k)
frame_vm_group_bin_7277 = frame (4k)
frame_vm_group_bin_7278 = frame (4k)
frame_vm_group_bin_7279 = frame (4k)
frame_vm_group_bin_7280 = frame (4k)
frame_vm_group_bin_7281 = frame (4k)
frame_vm_group_bin_7282 = frame (4k)
frame_vm_group_bin_7283 = frame (4k)
frame_vm_group_bin_7284 = frame (4k)
frame_vm_group_bin_7285 = frame (4k)
frame_vm_group_bin_7286 = frame (4k)
frame_vm_group_bin_7287 = frame (4k)
frame_vm_group_bin_7288 = frame (4k)
frame_vm_group_bin_7289 = frame (4k)
frame_vm_group_bin_7290 = frame (4k)
frame_vm_group_bin_7291 = frame (4k)
frame_vm_group_bin_7292 = frame (4k)
frame_vm_group_bin_7293 = frame (4k)
frame_vm_group_bin_7294 = frame (4k)
frame_vm_group_bin_7295 = frame (4k)
frame_vm_group_bin_7296 = frame (4k)
frame_vm_group_bin_7297 = frame (4k)
frame_vm_group_bin_7298 = frame (4k)
frame_vm_group_bin_7299 = frame (4k)
frame_vm_group_bin_7300 = frame (4k)
frame_vm_group_bin_7301 = frame (4k)
frame_vm_group_bin_7302 = frame (4k)
frame_vm_group_bin_7303 = frame (4k)
frame_vm_group_bin_7304 = frame (4k)
frame_vm_group_bin_7305 = frame (4k)
frame_vm_group_bin_7306 = frame (4k)
frame_vm_group_bin_7307 = frame (4k)
frame_vm_group_bin_7308 = frame (4k)
frame_vm_group_bin_7309 = frame (4k)
frame_vm_group_bin_7310 = frame (4k)
frame_vm_group_bin_7311 = frame (4k)
frame_vm_group_bin_7312 = frame (4k)
frame_vm_group_bin_7313 = frame (4k)
frame_vm_group_bin_7314 = frame (4k)
frame_vm_group_bin_7315 = frame (4k)
frame_vm_group_bin_7316 = frame (4k)
frame_vm_group_bin_7317 = frame (4k)
frame_vm_group_bin_7318 = frame (4k)
frame_vm_group_bin_7319 = frame (4k)
frame_vm_group_bin_7320 = frame (4k)
frame_vm_group_bin_7321 = frame (4k)
frame_vm_group_bin_7322 = frame (4k)
frame_vm_group_bin_7323 = frame (4k)
frame_vm_group_bin_7324 = frame (4k)
frame_vm_group_bin_7325 = frame (4k)
frame_vm_group_bin_7326 = frame (4k)
frame_vm_group_bin_7327 = frame (4k)
frame_vm_group_bin_7328 = frame (4k)
frame_vm_group_bin_7329 = frame (4k)
frame_vm_group_bin_7330 = frame (4k)
frame_vm_group_bin_7331 = frame (4k)
frame_vm_group_bin_7332 = frame (4k)
frame_vm_group_bin_7333 = frame (4k)
frame_vm_group_bin_7334 = frame (4k)
frame_vm_group_bin_7335 = frame (4k)
frame_vm_group_bin_7336 = frame (4k)
frame_vm_group_bin_7337 = frame (4k)
frame_vm_group_bin_7338 = frame (4k)
frame_vm_group_bin_7339 = frame (4k)
frame_vm_group_bin_7340 = frame (4k)
frame_vm_group_bin_7341 = frame (4k)
frame_vm_group_bin_7342 = frame (4k)
frame_vm_group_bin_7343 = frame (4k)
frame_vm_group_bin_7344 = frame (4k)
frame_vm_group_bin_7345 = frame (4k)
frame_vm_group_bin_7346 = frame (4k)
frame_vm_group_bin_7347 = frame (4k)
frame_vm_group_bin_7348 = frame (4k)
frame_vm_group_bin_7349 = frame (4k)
frame_vm_group_bin_7350 = frame (4k)
frame_vm_group_bin_7351 = frame (4k)
frame_vm_group_bin_7352 = frame (4k)
frame_vm_group_bin_7353 = frame (4k)
frame_vm_group_bin_7354 = frame (4k)
frame_vm_group_bin_7355 = frame (4k)
frame_vm_group_bin_7356 = frame (4k)
frame_vm_group_bin_7357 = frame (4k)
frame_vm_group_bin_7358 = frame (4k)
frame_vm_group_bin_7359 = frame (4k)
frame_vm_group_bin_7360 = frame (4k)
frame_vm_group_bin_7361 = frame (4k)
frame_vm_group_bin_7362 = frame (4k)
frame_vm_group_bin_7363 = frame (4k)
frame_vm_group_bin_7364 = frame (4k)
frame_vm_group_bin_7365 = frame (4k)
frame_vm_group_bin_7366 = frame (4k)
frame_vm_group_bin_7367 = frame (4k)
frame_vm_group_bin_7368 = frame (4k)
frame_vm_group_bin_7369 = frame (4k)
frame_vm_group_bin_7370 = frame (4k)
frame_vm_group_bin_7371 = frame (4k)
frame_vm_group_bin_7372 = frame (4k)
frame_vm_group_bin_7373 = frame (4k)
frame_vm_group_bin_7374 = frame (4k)
frame_vm_group_bin_7375 = frame (4k)
frame_vm_group_bin_7376 = frame (4k)
frame_vm_group_bin_7377 = frame (4k)
frame_vm_group_bin_7378 = frame (4k)
frame_vm_group_bin_7379 = frame (4k)
frame_vm_group_bin_7380 = frame (4k)
frame_vm_group_bin_7381 = frame (4k)
frame_vm_group_bin_7382 = frame (4k)
frame_vm_group_bin_7383 = frame (4k)
frame_vm_group_bin_7384 = frame (4k)
frame_vm_group_bin_7385 = frame (4k)
frame_vm_group_bin_7386 = frame (4k)
frame_vm_group_bin_7387 = frame (4k)
frame_vm_group_bin_7388 = frame (4k)
frame_vm_group_bin_7389 = frame (4k)
frame_vm_group_bin_7390 = frame (4k)
frame_vm_group_bin_7391 = frame (4k)
frame_vm_group_bin_7392 = frame (4k)
frame_vm_group_bin_7393 = frame (4k)
frame_vm_group_bin_7394 = frame (4k)
frame_vm_group_bin_7395 = frame (4k)
frame_vm_group_bin_7396 = frame (4k)
frame_vm_group_bin_7397 = frame (4k)
frame_vm_group_bin_7398 = frame (4k)
frame_vm_group_bin_7399 = frame (4k)
frame_vm_group_bin_7400 = frame (4k)
frame_vm_group_bin_7401 = frame (4k)
frame_vm_group_bin_7402 = frame (4k)
frame_vm_group_bin_7403 = frame (4k)
frame_vm_group_bin_7404 = frame (4k)
frame_vm_group_bin_7405 = frame (4k)
frame_vm_group_bin_7406 = frame (4k)
frame_vm_group_bin_7407 = frame (4k)
frame_vm_group_bin_7408 = frame (4k)
frame_vm_group_bin_7409 = frame (4k)
frame_vm_group_bin_7410 = frame (4k)
frame_vm_group_bin_7411 = frame (4k)
frame_vm_group_bin_7412 = frame (4k)
frame_vm_group_bin_7413 = frame (4k)
frame_vm_group_bin_7414 = frame (4k)
frame_vm_group_bin_7415 = frame (4k)
frame_vm_group_bin_7416 = frame (4k)
frame_vm_group_bin_7417 = frame (4k)
frame_vm_group_bin_7418 = frame (4k)
frame_vm_group_bin_7419 = frame (4k)
frame_vm_group_bin_7420 = frame (4k)
frame_vm_group_bin_7421 = frame (4k)
frame_vm_group_bin_7422 = frame (4k)
frame_vm_group_bin_7423 = frame (4k)
frame_vm_group_bin_7424 = frame (4k)
frame_vm_group_bin_7425 = frame (4k)
frame_vm_group_bin_7426 = frame (4k)
frame_vm_group_bin_7427 = frame (4k)
frame_vm_group_bin_7428 = frame (4k)
frame_vm_group_bin_7429 = frame (4k)
frame_vm_group_bin_7430 = frame (4k)
frame_vm_group_bin_7431 = frame (4k)
frame_vm_group_bin_7432 = frame (4k)
frame_vm_group_bin_7433 = frame (4k)
frame_vm_group_bin_7434 = frame (4k)
frame_vm_group_bin_7435 = frame (4k)
frame_vm_group_bin_7436 = frame (4k)
frame_vm_group_bin_7437 = frame (4k)
frame_vm_group_bin_7438 = frame (4k)
frame_vm_group_bin_7439 = frame (4k)
frame_vm_group_bin_7440 = frame (4k)
frame_vm_group_bin_7441 = frame (4k)
frame_vm_group_bin_7442 = frame (4k)
frame_vm_group_bin_7443 = frame (4k)
frame_vm_group_bin_7444 = frame (4k)
frame_vm_group_bin_7445 = frame (4k)
frame_vm_group_bin_7446 = frame (4k)
frame_vm_group_bin_7447 = frame (4k)
frame_vm_group_bin_7448 = frame (4k)
frame_vm_group_bin_7449 = frame (4k)
frame_vm_group_bin_7450 = frame (4k)
frame_vm_group_bin_7451 = frame (4k)
frame_vm_group_bin_7452 = frame (4k)
frame_vm_group_bin_7453 = frame (4k)
frame_vm_group_bin_7454 = frame (4k)
frame_vm_group_bin_7455 = frame (4k)
frame_vm_group_bin_7456 = frame (4k)
frame_vm_group_bin_7457 = frame (4k)
frame_vm_group_bin_7458 = frame (4k)
frame_vm_group_bin_7459 = frame (4k)
frame_vm_group_bin_7460 = frame (4k)
frame_vm_group_bin_7461 = frame (4k)
frame_vm_group_bin_7462 = frame (4k)
frame_vm_group_bin_7463 = frame (4k)
frame_vm_group_bin_7464 = frame (4k)
frame_vm_group_bin_7465 = frame (4k)
frame_vm_group_bin_7466 = frame (4k)
frame_vm_group_bin_7467 = frame (4k)
frame_vm_group_bin_7468 = frame (4k)
frame_vm_group_bin_7469 = frame (4k)
frame_vm_group_bin_7470 = frame (4k)
frame_vm_group_bin_7471 = frame (4k)
frame_vm_group_bin_7472 = frame (4k)
frame_vm_group_bin_7473 = frame (4k)
frame_vm_group_bin_7474 = frame (4k)
frame_vm_group_bin_7475 = frame (4k)
frame_vm_group_bin_7476 = frame (4k)
frame_vm_group_bin_7477 = frame (4k)
frame_vm_group_bin_7478 = frame (4k)
frame_vm_group_bin_7479 = frame (4k)
frame_vm_group_bin_7480 = frame (4k)
frame_vm_group_bin_7481 = frame (4k)
frame_vm_group_bin_7482 = frame (4k)
frame_vm_group_bin_7483 = frame (4k)
frame_vm_group_bin_7484 = frame (4k)
frame_vm_group_bin_7485 = frame (4k)
frame_vm_group_bin_7486 = frame (4k)
frame_vm_group_bin_7487 = frame (4k)
frame_vm_group_bin_7488 = frame (4k)
frame_vm_group_bin_7489 = frame (4k)
frame_vm_group_bin_7490 = frame (4k)
frame_vm_group_bin_7491 = frame (4k)
frame_vm_group_bin_7492 = frame (4k)
frame_vm_group_bin_7493 = frame (4k)
frame_vm_group_bin_7494 = frame (4k)
frame_vm_group_bin_7495 = frame (4k)
frame_vm_group_bin_7496 = frame (4k)
frame_vm_group_bin_7497 = frame (4k)
frame_vm_group_bin_7498 = frame (4k)
frame_vm_group_bin_7499 = frame (4k)
frame_vm_group_bin_7500 = frame (4k)
frame_vm_group_bin_7501 = frame (4k)
frame_vm_group_bin_7502 = frame (4k)
frame_vm_group_bin_7503 = frame (4k)
frame_vm_group_bin_7504 = frame (4k)
frame_vm_group_bin_7505 = frame (4k)
frame_vm_group_bin_7506 = frame (4k)
frame_vm_group_bin_7507 = frame (4k)
frame_vm_group_bin_7508 = frame (4k)
frame_vm_group_bin_7509 = frame (4k)
frame_vm_group_bin_7510 = frame (4k)
frame_vm_group_bin_7511 = frame (4k)
frame_vm_group_bin_7512 = frame (4k)
frame_vm_group_bin_7513 = frame (4k)
frame_vm_group_bin_7514 = frame (4k)
frame_vm_group_bin_7515 = frame (4k)
frame_vm_group_bin_7516 = frame (4k)
frame_vm_group_bin_7517 = frame (4k)
frame_vm_group_bin_7518 = frame (4k)
frame_vm_group_bin_7519 = frame (4k)
frame_vm_group_bin_7520 = frame (4k)
frame_vm_group_bin_7521 = frame (4k)
frame_vm_group_bin_7522 = frame (4k)
frame_vm_group_bin_7523 = frame (4k)
frame_vm_group_bin_7524 = frame (4k)
frame_vm_group_bin_7525 = frame (4k)
frame_vm_group_bin_7526 = frame (4k)
frame_vm_group_bin_7527 = frame (4k)
frame_vm_group_bin_7528 = frame (4k)
frame_vm_group_bin_7529 = frame (4k)
frame_vm_group_bin_7530 = frame (4k)
frame_vm_group_bin_7531 = frame (4k)
frame_vm_group_bin_7532 = frame (4k)
frame_vm_group_bin_7533 = frame (4k)
frame_vm_group_bin_7534 = frame (4k)
frame_vm_group_bin_7535 = frame (4k)
frame_vm_group_bin_7536 = frame (4k)
frame_vm_group_bin_7537 = frame (4k)
frame_vm_group_bin_7538 = frame (4k)
frame_vm_group_bin_7539 = frame (4k)
frame_vm_group_bin_7540 = frame (4k)
frame_vm_group_bin_7541 = frame (4k)
frame_vm_group_bin_7542 = frame (4k)
frame_vm_group_bin_7543 = frame (4k)
frame_vm_group_bin_7544 = frame (4k)
frame_vm_group_bin_7545 = frame (4k)
frame_vm_group_bin_7546 = frame (4k)
frame_vm_group_bin_7547 = frame (4k)
frame_vm_group_bin_7548 = frame (4k)
frame_vm_group_bin_7549 = frame (4k)
frame_vm_group_bin_7550 = frame (4k)
frame_vm_group_bin_7551 = frame (4k)
frame_vm_group_bin_7552 = frame (4k)
frame_vm_group_bin_7553 = frame (4k)
frame_vm_group_bin_7554 = frame (4k)
frame_vm_group_bin_7555 = frame (4k)
frame_vm_group_bin_7556 = frame (4k)
frame_vm_group_bin_7557 = frame (4k)
frame_vm_group_bin_7558 = frame (4k)
frame_vm_group_bin_7559 = frame (4k)
frame_vm_group_bin_7560 = frame (4k)
frame_vm_group_bin_7561 = frame (4k)
frame_vm_group_bin_7562 = frame (4k)
frame_vm_group_bin_7563 = frame (4k)
frame_vm_group_bin_7564 = frame (4k)
frame_vm_group_bin_7565 = frame (4k)
frame_vm_group_bin_7566 = frame (4k)
frame_vm_group_bin_7567 = frame (4k)
frame_vm_group_bin_7568 = frame (4k)
frame_vm_group_bin_7569 = frame (4k)
frame_vm_group_bin_7570 = frame (4k)
frame_vm_group_bin_7571 = frame (4k)
frame_vm_group_bin_7572 = frame (4k)
frame_vm_group_bin_7573 = frame (4k)
frame_vm_group_bin_7574 = frame (4k)
frame_vm_group_bin_7575 = frame (4k)
frame_vm_group_bin_7576 = frame (4k)
frame_vm_group_bin_7577 = frame (4k)
frame_vm_group_bin_7578 = frame (4k)
frame_vm_group_bin_7579 = frame (4k)
frame_vm_group_bin_7580 = frame (4k)
frame_vm_group_bin_7581 = frame (4k)
frame_vm_group_bin_7582 = frame (4k)
frame_vm_group_bin_7583 = frame (4k)
frame_vm_group_bin_7584 = frame (4k)
frame_vm_group_bin_7585 = frame (4k)
frame_vm_group_bin_7586 = frame (4k)
frame_vm_group_bin_7587 = frame (4k)
frame_vm_group_bin_7588 = frame (4k)
frame_vm_group_bin_7589 = frame (4k)
frame_vm_group_bin_7590 = frame (4k)
frame_vm_group_bin_7591 = frame (4k)
frame_vm_group_bin_7592 = frame (4k)
frame_vm_group_bin_7593 = frame (4k)
frame_vm_group_bin_7594 = frame (4k)
frame_vm_group_bin_7595 = frame (4k)
frame_vm_group_bin_7596 = frame (4k)
frame_vm_group_bin_7597 = frame (4k)
frame_vm_group_bin_7598 = frame (4k)
frame_vm_group_bin_7599 = frame (4k)
frame_vm_group_bin_7600 = frame (4k)
frame_vm_group_bin_7601 = frame (4k)
frame_vm_group_bin_7602 = frame (4k)
frame_vm_group_bin_7603 = frame (4k)
frame_vm_group_bin_7604 = frame (4k)
frame_vm_group_bin_7605 = frame (4k)
frame_vm_group_bin_7606 = frame (4k)
frame_vm_group_bin_7607 = frame (4k)
frame_vm_group_bin_7608 = frame (4k)
frame_vm_group_bin_7609 = frame (4k)
frame_vm_group_bin_7610 = frame (4k)
frame_vm_group_bin_7611 = frame (4k)
frame_vm_group_bin_7612 = frame (4k)
frame_vm_group_bin_7613 = frame (4k)
frame_vm_group_bin_7614 = frame (4k)
frame_vm_group_bin_7615 = frame (4k)
frame_vm_group_bin_7616 = frame (4k)
frame_vm_group_bin_7617 = frame (4k)
frame_vm_group_bin_7618 = frame (4k)
frame_vm_group_bin_7619 = frame (4k)
frame_vm_group_bin_7620 = frame (4k)
frame_vm_group_bin_7621 = frame (4k)
frame_vm_group_bin_7622 = frame (4k)
frame_vm_group_bin_7623 = frame (4k)
frame_vm_group_bin_7624 = frame (4k)
frame_vm_group_bin_7625 = frame (4k)
frame_vm_group_bin_7626 = frame (4k)
frame_vm_group_bin_7627 = frame (4k)
frame_vm_group_bin_7628 = frame (4k)
frame_vm_group_bin_7629 = frame (4k)
frame_vm_group_bin_7630 = frame (4k)
frame_vm_group_bin_7631 = frame (4k)
frame_vm_group_bin_7632 = frame (4k)
frame_vm_group_bin_7633 = frame (4k)
frame_vm_group_bin_7634 = frame (4k)
frame_vm_group_bin_7635 = frame (4k)
frame_vm_group_bin_7636 = frame (4k)
frame_vm_group_bin_7637 = frame (4k)
frame_vm_group_bin_7638 = frame (4k)
frame_vm_group_bin_7639 = frame (4k)
frame_vm_group_bin_7640 = frame (4k)
frame_vm_group_bin_7641 = frame (4k)
frame_vm_group_bin_7642 = frame (4k)
frame_vm_group_bin_7643 = frame (4k)
frame_vm_group_bin_7644 = frame (4k)
frame_vm_group_bin_7645 = frame (4k)
frame_vm_group_bin_7646 = frame (4k)
frame_vm_group_bin_7647 = frame (4k)
frame_vm_group_bin_7648 = frame (4k)
frame_vm_group_bin_7649 = frame (4k)
frame_vm_group_bin_7650 = frame (4k)
frame_vm_group_bin_7651 = frame (4k)
frame_vm_group_bin_7652 = frame (4k)
frame_vm_group_bin_7653 = frame (4k)
frame_vm_group_bin_7654 = frame (4k)
frame_vm_group_bin_7655 = frame (4k)
frame_vm_group_bin_7656 = frame (4k)
frame_vm_group_bin_7657 = frame (4k)
frame_vm_group_bin_7658 = frame (4k)
frame_vm_group_bin_7659 = frame (4k)
frame_vm_group_bin_7660 = frame (4k)
frame_vm_group_bin_7661 = frame (4k)
frame_vm_group_bin_7662 = frame (4k)
frame_vm_group_bin_7663 = frame (4k)
frame_vm_group_bin_7664 = frame (4k)
frame_vm_group_bin_7665 = frame (4k)
frame_vm_group_bin_7666 = frame (4k)
frame_vm_group_bin_7667 = frame (4k)
frame_vm_group_bin_7668 = frame (4k)
frame_vm_group_bin_7669 = frame (4k)
frame_vm_group_bin_7670 = frame (4k)
frame_vm_group_bin_7671 = frame (4k)
frame_vm_group_bin_7672 = frame (4k)
frame_vm_group_bin_7673 = frame (4k)
frame_vm_group_bin_7674 = frame (4k)
frame_vm_group_bin_7675 = frame (4k)
frame_vm_group_bin_7676 = frame (4k)
frame_vm_group_bin_7677 = frame (4k)
frame_vm_group_bin_7678 = frame (4k)
frame_vm_group_bin_7679 = frame (4k)
frame_vm_group_bin_7680 = frame (4k)
frame_vm_group_bin_7681 = frame (4k)
frame_vm_group_bin_7682 = frame (4k)
frame_vm_group_bin_7683 = frame (4k)
frame_vm_group_bin_7684 = frame (4k)
frame_vm_group_bin_7685 = frame (4k)
frame_vm_group_bin_7686 = frame (4k)
frame_vm_group_bin_7687 = frame (4k)
frame_vm_group_bin_7688 = frame (4k)
frame_vm_group_bin_7689 = frame (4k)
frame_vm_group_bin_7690 = frame (4k)
frame_vm_group_bin_7691 = frame (4k)
frame_vm_group_bin_7692 = frame (4k)
frame_vm_group_bin_7693 = frame (4k)
frame_vm_group_bin_7694 = frame (4k)
frame_vm_group_bin_7695 = frame (4k)
frame_vm_group_bin_7696 = frame (4k)
frame_vm_group_bin_7697 = frame (4k)
frame_vm_group_bin_7698 = frame (4k)
frame_vm_group_bin_7699 = frame (4k)
frame_vm_group_bin_7700 = frame (4k)
frame_vm_group_bin_7701 = frame (4k)
frame_vm_group_bin_7702 = frame (4k)
frame_vm_group_bin_7703 = frame (4k)
frame_vm_group_bin_7704 = frame (4k)
frame_vm_group_bin_7705 = frame (4k)
frame_vm_group_bin_7706 = frame (4k)
frame_vm_group_bin_7707 = frame (4k)
frame_vm_group_bin_7708 = frame (4k)
frame_vm_group_bin_7709 = frame (4k)
frame_vm_group_bin_7710 = frame (4k)
frame_vm_group_bin_7711 = frame (4k)
frame_vm_group_bin_7712 = frame (4k)
frame_vm_group_bin_7713 = frame (4k)
frame_vm_group_bin_7714 = frame (4k)
frame_vm_group_bin_7715 = frame (4k)
frame_vm_group_bin_7716 = frame (4k)
frame_vm_group_bin_7717 = frame (4k)
frame_vm_group_bin_7718 = frame (4k)
frame_vm_group_bin_7719 = frame (4k)
frame_vm_group_bin_7720 = frame (4k)
frame_vm_group_bin_7721 = frame (4k)
frame_vm_group_bin_7722 = frame (4k)
frame_vm_group_bin_7723 = frame (4k)
frame_vm_group_bin_7724 = frame (4k)
frame_vm_group_bin_7725 = frame (4k)
frame_vm_group_bin_7726 = frame (4k)
frame_vm_group_bin_7727 = frame (4k)
frame_vm_group_bin_7728 = frame (4k)
frame_vm_group_bin_7729 = frame (4k)
frame_vm_group_bin_7730 = frame (4k)
frame_vm_group_bin_7731 = frame (4k)
frame_vm_group_bin_7732 = frame (4k)
frame_vm_group_bin_7733 = frame (4k)
frame_vm_group_bin_7734 = frame (4k)
frame_vm_group_bin_7735 = frame (4k)
frame_vm_group_bin_7736 = frame (4k)
frame_vm_group_bin_7737 = frame (4k)
frame_vm_group_bin_7738 = frame (4k)
frame_vm_group_bin_7739 = frame (4k)
frame_vm_group_bin_7740 = frame (4k)
frame_vm_group_bin_7741 = frame (4k)
frame_vm_group_bin_7742 = frame (4k)
frame_vm_group_bin_7743 = frame (4k)
frame_vm_group_bin_7744 = frame (4k)
frame_vm_group_bin_7745 = frame (4k)
frame_vm_group_bin_7746 = frame (4k)
frame_vm_group_bin_7747 = frame (4k)
frame_vm_group_bin_7748 = frame (4k)
frame_vm_group_bin_7749 = frame (4k)
frame_vm_group_bin_7750 = frame (4k)
frame_vm_group_bin_7751 = frame (4k)
frame_vm_group_bin_7752 = frame (4k)
frame_vm_group_bin_7753 = frame (4k)
frame_vm_group_bin_7754 = frame (4k)
frame_vm_group_bin_7755 = frame (4k)
frame_vm_group_bin_7756 = frame (4k)
frame_vm_group_bin_7757 = frame (4k)
frame_vm_group_bin_7758 = frame (4k)
frame_vm_group_bin_7759 = frame (4k)
frame_vm_group_bin_7760 = frame (4k)
frame_vm_group_bin_7761 = frame (4k)
frame_vm_group_bin_7762 = frame (4k)
frame_vm_group_bin_7763 = frame (4k)
frame_vm_group_bin_7764 = frame (4k)
frame_vm_group_bin_7765 = frame (4k)
frame_vm_group_bin_7766 = frame (4k)
frame_vm_group_bin_7767 = frame (4k)
frame_vm_group_bin_7768 = frame (4k)
frame_vm_group_bin_7769 = frame (4k)
frame_vm_group_bin_7770 = frame (4k)
frame_vm_group_bin_7771 = frame (4k)
frame_vm_group_bin_7772 = frame (4k)
frame_vm_group_bin_7773 = frame (4k)
frame_vm_group_bin_7774 = frame (4k)
frame_vm_group_bin_7775 = frame (4k)
frame_vm_group_bin_7776 = frame (4k)
frame_vm_group_bin_7777 = frame (4k)
frame_vm_group_bin_7778 = frame (4k)
frame_vm_group_bin_7779 = frame (4k)
frame_vm_group_bin_7780 = frame (4k)
frame_vm_group_bin_7781 = frame (4k)
frame_vm_group_bin_7782 = frame (4k)
frame_vm_group_bin_7783 = frame (4k)
frame_vm_group_bin_7784 = frame (4k)
frame_vm_group_bin_7785 = frame (4k)
frame_vm_group_bin_7786 = frame (4k)
frame_vm_group_bin_7787 = frame (4k)
frame_vm_group_bin_7788 = frame (4k)
frame_vm_group_bin_7789 = frame (4k)
frame_vm_group_bin_7790 = frame (4k)
frame_vm_group_bin_7791 = frame (4k)
frame_vm_group_bin_7792 = frame (4k)
frame_vm_group_bin_7793 = frame (4k)
frame_vm_group_bin_7794 = frame (4k)
frame_vm_group_bin_7795 = frame (4k)
frame_vm_group_bin_7796 = frame (4k)
frame_vm_group_bin_7797 = frame (4k)
frame_vm_group_bin_7798 = frame (4k)
frame_vm_group_bin_7799 = frame (4k)
frame_vm_group_bin_7800 = frame (4k)
frame_vm_group_bin_7801 = frame (4k)
frame_vm_group_bin_7802 = frame (4k)
frame_vm_group_bin_7803 = frame (4k)
frame_vm_group_bin_7804 = frame (4k)
frame_vm_group_bin_7805 = frame (4k)
frame_vm_group_bin_7806 = frame (4k)
frame_vm_group_bin_7807 = frame (4k)
frame_vm_group_bin_7808 = frame (4k)
frame_vm_group_bin_7809 = frame (4k)
frame_vm_group_bin_7810 = frame (4k)
frame_vm_group_bin_7811 = frame (4k)
frame_vm_group_bin_7812 = frame (4k)
frame_vm_group_bin_7813 = frame (4k)
frame_vm_group_bin_7814 = frame (4k)
frame_vm_group_bin_7815 = frame (4k)
frame_vm_group_bin_7816 = frame (4k)
frame_vm_group_bin_7817 = frame (4k)
frame_vm_group_bin_7818 = frame (4k)
frame_vm_group_bin_7819 = frame (4k)
frame_vm_group_bin_7820 = frame (4k)
frame_vm_group_bin_7821 = frame (4k)
frame_vm_group_bin_7822 = frame (4k)
frame_vm_group_bin_7823 = frame (4k)
frame_vm_group_bin_7824 = frame (4k)
frame_vm_group_bin_7825 = frame (4k)
frame_vm_group_bin_7826 = frame (4k)
frame_vm_group_bin_7827 = frame (4k)
frame_vm_group_bin_7828 = frame (4k)
frame_vm_group_bin_7829 = frame (4k)
frame_vm_group_bin_7830 = frame (4k)
frame_vm_group_bin_7831 = frame (4k)
frame_vm_group_bin_7832 = frame (4k)
frame_vm_group_bin_7833 = frame (4k)
frame_vm_group_bin_7834 = frame (4k)
frame_vm_group_bin_7835 = frame (4k)
frame_vm_group_bin_7836 = frame (4k)
frame_vm_group_bin_7837 = frame (4k)
frame_vm_group_bin_7838 = frame (4k)
frame_vm_group_bin_7839 = frame (4k)
frame_vm_group_bin_7840 = frame (4k)
frame_vm_group_bin_7841 = frame (4k)
frame_vm_group_bin_7842 = frame (4k)
frame_vm_group_bin_7843 = frame (4k)
frame_vm_group_bin_7844 = frame (4k)
frame_vm_group_bin_7845 = frame (4k)
frame_vm_group_bin_7846 = frame (4k)
frame_vm_group_bin_7847 = frame (4k)
frame_vm_group_bin_7848 = frame (4k)
frame_vm_group_bin_7849 = frame (4k)
frame_vm_group_bin_7850 = frame (4k)
frame_vm_group_bin_7851 = frame (4k)
frame_vm_group_bin_7852 = frame (4k)
frame_vm_group_bin_7853 = frame (4k)
frame_vm_group_bin_7854 = frame (4k)
frame_vm_group_bin_7855 = frame (4k)
frame_vm_group_bin_7856 = frame (4k)
frame_vm_group_bin_7857 = frame (4k)
frame_vm_group_bin_7858 = frame (4k)
frame_vm_group_bin_7859 = frame (4k)
frame_vm_group_bin_7860 = frame (4k)
frame_vm_group_bin_7861 = frame (4k)
frame_vm_group_bin_7862 = frame (4k)
frame_vm_group_bin_7863 = frame (4k)
frame_vm_group_bin_7864 = frame (4k)
frame_vm_group_bin_7865 = frame (4k)
frame_vm_group_bin_7866 = frame (4k)
frame_vm_group_bin_7867 = frame (4k)
frame_vm_group_bin_7868 = frame (4k)
frame_vm_group_bin_7869 = frame (4k)
frame_vm_group_bin_7870 = frame (4k)
frame_vm_group_bin_7871 = frame (4k)
frame_vm_group_bin_7872 = frame (4k)
frame_vm_group_bin_7873 = frame (4k)
frame_vm_group_bin_7874 = frame (4k)
frame_vm_group_bin_7875 = frame (4k)
frame_vm_group_bin_7876 = frame (4k)
frame_vm_group_bin_7877 = frame (4k)
frame_vm_group_bin_7878 = frame (4k)
frame_vm_group_bin_7879 = frame (4k)
frame_vm_group_bin_7880 = frame (4k)
frame_vm_group_bin_7881 = frame (4k)
frame_vm_group_bin_7882 = frame (4k)
frame_vm_group_bin_7883 = frame (4k)
frame_vm_group_bin_7884 = frame (4k)
frame_vm_group_bin_7885 = frame (4k)
frame_vm_group_bin_7886 = frame (4k)
frame_vm_group_bin_7887 = frame (4k)
frame_vm_group_bin_7888 = frame (4k)
frame_vm_group_bin_7889 = frame (4k)
frame_vm_group_bin_7890 = frame (4k)
frame_vm_group_bin_7891 = frame (4k)
frame_vm_group_bin_7892 = frame (4k)
frame_vm_group_bin_7893 = frame (4k)
frame_vm_group_bin_7894 = frame (4k)
frame_vm_group_bin_7895 = frame (4k)
frame_vm_group_bin_7896 = frame (4k)
frame_vm_group_bin_7897 = frame (4k)
frame_vm_group_bin_7898 = frame (4k)
frame_vm_group_bin_7899 = frame (4k)
frame_vm_group_bin_7900 = frame (4k)
frame_vm_group_bin_7901 = frame (4k)
frame_vm_group_bin_7902 = frame (4k)
frame_vm_group_bin_7903 = frame (4k)
frame_vm_group_bin_7904 = frame (4k)
frame_vm_group_bin_7905 = frame (4k)
frame_vm_group_bin_7906 = frame (4k)
frame_vm_group_bin_7907 = frame (4k)
frame_vm_group_bin_7908 = frame (4k)
frame_vm_group_bin_7909 = frame (4k)
frame_vm_group_bin_7910 = frame (4k)
frame_vm_group_bin_7911 = frame (4k)
frame_vm_group_bin_7912 = frame (4k)
frame_vm_group_bin_7913 = frame (4k)
frame_vm_group_bin_7914 = frame (4k)
frame_vm_group_bin_7915 = frame (4k)
frame_vm_group_bin_7916 = frame (4k)
frame_vm_group_bin_7917 = frame (4k)
frame_vm_group_bin_7918 = frame (4k)
frame_vm_group_bin_7919 = frame (4k)
frame_vm_group_bin_7920 = frame (4k)
frame_vm_group_bin_7921 = frame (4k)
frame_vm_group_bin_7922 = frame (4k)
frame_vm_group_bin_7923 = frame (4k)
frame_vm_group_bin_7924 = frame (4k)
frame_vm_group_bin_7925 = frame (4k)
frame_vm_group_bin_7926 = frame (4k)
frame_vm_group_bin_7927 = frame (4k)
frame_vm_group_bin_7928 = frame (4k)
frame_vm_group_bin_7929 = frame (4k)
frame_vm_group_bin_7930 = frame (4k)
frame_vm_group_bin_7931 = frame (4k)
frame_vm_group_bin_7932 = frame (4k)
frame_vm_group_bin_7933 = frame (4k)
frame_vm_group_bin_7934 = frame (4k)
frame_vm_group_bin_7935 = frame (4k)
frame_vm_group_bin_7936 = frame (4k)
frame_vm_group_bin_7937 = frame (4k)
frame_vm_group_bin_7938 = frame (4k)
frame_vm_group_bin_7939 = frame (4k)
frame_vm_group_bin_7940 = frame (4k)
frame_vm_group_bin_7941 = frame (4k)
frame_vm_group_bin_7942 = frame (4k)
frame_vm_group_bin_7943 = frame (4k)
frame_vm_group_bin_7944 = frame (4k)
frame_vm_group_bin_7945 = frame (4k)
frame_vm_group_bin_7946 = frame (4k)
frame_vm_group_bin_7947 = frame (4k)
frame_vm_group_bin_7948 = frame (4k)
frame_vm_group_bin_7949 = frame (4k)
frame_vm_group_bin_7950 = frame (4k)
frame_vm_group_bin_7951 = frame (4k)
frame_vm_group_bin_7952 = frame (4k)
frame_vm_group_bin_7953 = frame (4k)
frame_vm_group_bin_7954 = frame (4k)
frame_vm_group_bin_7955 = frame (4k)
frame_vm_group_bin_7956 = frame (4k)
frame_vm_group_bin_7957 = frame (4k)
frame_vm_group_bin_7958 = frame (4k)
frame_vm_group_bin_7959 = frame (4k)
frame_vm_group_bin_7960 = frame (4k)
frame_vm_group_bin_7961 = frame (4k)
frame_vm_group_bin_7962 = frame (4k)
frame_vm_group_bin_7963 = frame (4k)
frame_vm_group_bin_7964 = frame (4k)
frame_vm_group_bin_7965 = frame (4k)
frame_vm_group_bin_7966 = frame (4k)
frame_vm_group_bin_7967 = frame (4k)
frame_vm_group_bin_7968 = frame (4k)
frame_vm_group_bin_7969 = frame (4k)
frame_vm_group_bin_7970 = frame (4k)
frame_vm_group_bin_7971 = frame (4k)
frame_vm_group_bin_7972 = frame (4k)
frame_vm_group_bin_7973 = frame (4k)
frame_vm_group_bin_7974 = frame (4k)
frame_vm_group_bin_7975 = frame (4k)
frame_vm_group_bin_7976 = frame (4k)
frame_vm_group_bin_7977 = frame (4k)
frame_vm_group_bin_7978 = frame (4k)
frame_vm_group_bin_7979 = frame (4k)
frame_vm_group_bin_7980 = frame (4k)
frame_vm_group_bin_7981 = frame (4k)
frame_vm_group_bin_7982 = frame (4k)
frame_vm_group_bin_7983 = frame (4k)
frame_vm_group_bin_7984 = frame (4k)
frame_vm_group_bin_7985 = frame (4k)
frame_vm_group_bin_7986 = frame (4k)
frame_vm_group_bin_7987 = frame (4k)
frame_vm_group_bin_7988 = frame (4k)
frame_vm_group_bin_7989 = frame (4k)
frame_vm_group_bin_7990 = frame (4k)
frame_vm_group_bin_7991 = frame (4k)
frame_vm_group_bin_7992 = frame (4k)
frame_vm_group_bin_7993 = frame (4k)
frame_vm_group_bin_7994 = frame (4k)
frame_vm_group_bin_7995 = frame (4k)
frame_vm_group_bin_7996 = frame (4k)
frame_vm_group_bin_7997 = frame (4k)
frame_vm_group_bin_7998 = frame (4k)
frame_vm_group_bin_7999 = frame (4k)
frame_vm_group_bin_8000 = frame (4k)
frame_vm_group_bin_8001 = frame (4k)
frame_vm_group_bin_8002 = frame (4k)
frame_vm_group_bin_8003 = frame (4k)
frame_vm_group_bin_8004 = frame (4k)
frame_vm_group_bin_8005 = frame (4k)
frame_vm_group_bin_8006 = frame (4k)
frame_vm_group_bin_8007 = frame (4k)
frame_vm_group_bin_8008 = frame (4k)
frame_vm_group_bin_8009 = frame (4k)
frame_vm_group_bin_8010 = frame (4k)
frame_vm_group_bin_8011 = frame (4k)
frame_vm_group_bin_8012 = frame (4k)
frame_vm_group_bin_8013 = frame (4k)
frame_vm_group_bin_8014 = frame (4k)
frame_vm_group_bin_8015 = frame (4k)
frame_vm_group_bin_8016 = frame (4k)
frame_vm_group_bin_8017 = frame (4k)
frame_vm_group_bin_8018 = frame (4k)
frame_vm_group_bin_8019 = frame (4k)
frame_vm_group_bin_8020 = frame (4k)
frame_vm_group_bin_8021 = frame (4k)
frame_vm_group_bin_8022 = frame (4k)
frame_vm_group_bin_8023 = frame (4k)
frame_vm_group_bin_8024 = frame (4k)
frame_vm_group_bin_8025 = frame (4k)
frame_vm_group_bin_8026 = frame (4k)
frame_vm_group_bin_8027 = frame (4k)
frame_vm_group_bin_8028 = frame (4k)
frame_vm_group_bin_8029 = frame (4k)
frame_vm_group_bin_8030 = frame (4k)
frame_vm_group_bin_8031 = frame (4k)
frame_vm_group_bin_8032 = frame (4k)
frame_vm_group_bin_8033 = frame (4k)
frame_vm_group_bin_8034 = frame (4k)
frame_vm_group_bin_8035 = frame (4k)
frame_vm_group_bin_8036 = frame (4k)
frame_vm_group_bin_8037 = frame (4k)
frame_vm_group_bin_8038 = frame (4k)
frame_vm_group_bin_8039 = frame (4k)
frame_vm_group_bin_8040 = frame (4k)
frame_vm_group_bin_8041 = frame (4k)
frame_vm_group_bin_8042 = frame (4k)
frame_vm_group_bin_8043 = frame (4k)
frame_vm_group_bin_8044 = frame (4k)
frame_vm_group_bin_8045 = frame (4k)
frame_vm_group_bin_8046 = frame (4k)
frame_vm_group_bin_8047 = frame (4k)
frame_vm_group_bin_8048 = frame (4k)
frame_vm_group_bin_8049 = frame (4k)
frame_vm_group_bin_8050 = frame (4k)
frame_vm_group_bin_8051 = frame (4k)
frame_vm_group_bin_8052 = frame (4k)
frame_vm_group_bin_8053 = frame (4k)
frame_vm_group_bin_8054 = frame (4k)
frame_vm_group_bin_8055 = frame (4k)
frame_vm_group_bin_8056 = frame (4k)
frame_vm_group_bin_8057 = frame (4k)
frame_vm_group_bin_8058 = frame (4k)
frame_vm_group_bin_8059 = frame (4k)
frame_vm_group_bin_8060 = frame (4k)
frame_vm_group_bin_8061 = frame (4k)
frame_vm_group_bin_8062 = frame (4k)
frame_vm_group_bin_8063 = frame (4k)
frame_vm_group_bin_8064 = frame (4k)
frame_vm_group_bin_8065 = frame (4k)
frame_vm_group_bin_8066 = frame (4k)
frame_vm_group_bin_8067 = frame (4k)
frame_vm_group_bin_8068 = frame (4k)
frame_vm_group_bin_8069 = frame (4k)
frame_vm_group_bin_8070 = frame (4k)
frame_vm_group_bin_8071 = frame (4k)
frame_vm_group_bin_8072 = frame (4k)
frame_vm_group_bin_8073 = frame (4k)
frame_vm_group_bin_8074 = frame (4k)
frame_vm_group_bin_8075 = frame (4k)
frame_vm_group_bin_8076 = frame (4k)
frame_vm_group_bin_8077 = frame (4k)
frame_vm_group_bin_8078 = frame (4k)
frame_vm_group_bin_8079 = frame (4k)
frame_vm_group_bin_8080 = frame (4k)
frame_vm_group_bin_8081 = frame (4k)
frame_vm_group_bin_8082 = frame (4k)
frame_vm_group_bin_8083 = frame (4k)
frame_vm_group_bin_8084 = frame (4k)
frame_vm_group_bin_8085 = frame (4k)
frame_vm_group_bin_8086 = frame (4k)
frame_vm_group_bin_8087 = frame (4k)
frame_vm_group_bin_8088 = frame (4k)
frame_vm_group_bin_8089 = frame (4k)
frame_vm_group_bin_8090 = frame (4k)
frame_vm_group_bin_8091 = frame (4k)
frame_vm_group_bin_8092 = frame (4k)
frame_vm_group_bin_8093 = frame (4k)
frame_vm_group_bin_8094 = frame (4k)
frame_vm_group_bin_8095 = frame (4k)
frame_vm_group_bin_8096 = frame (4k)
frame_vm_group_bin_8097 = frame (4k)
frame_vm_group_bin_8098 = frame (4k)
frame_vm_group_bin_8099 = frame (4k)
frame_vm_group_bin_8100 = frame (4k)
frame_vm_group_bin_8101 = frame (4k)
frame_vm_group_bin_8102 = frame (4k)
frame_vm_group_bin_8103 = frame (4k)
frame_vm_group_bin_8104 = frame (4k)
frame_vm_group_bin_8105 = frame (4k)
frame_vm_group_bin_8106 = frame (4k)
frame_vm_group_bin_8107 = frame (4k)
frame_vm_group_bin_8108 = frame (4k)
frame_vm_group_bin_8109 = frame (4k)
frame_vm_group_bin_8110 = frame (4k)
frame_vm_group_bin_8111 = frame (4k)
frame_vm_group_bin_8112 = frame (4k)
frame_vm_group_bin_8113 = frame (4k)
frame_vm_group_bin_8114 = frame (4k)
frame_vm_group_bin_8115 = frame (4k)
frame_vm_group_bin_8116 = frame (4k)
frame_vm_group_bin_8117 = frame (4k)
frame_vm_group_bin_8118 = frame (4k)
frame_vm_group_bin_8119 = frame (4k)
frame_vm_group_bin_8120 = frame (4k)
frame_vm_group_bin_8121 = frame (4k)
frame_vm_group_bin_8122 = frame (4k)
frame_vm_group_bin_8123 = frame (4k)
frame_vm_group_bin_8124 = frame (4k)
frame_vm_group_bin_8125 = frame (4k)
frame_vm_group_bin_8126 = frame (4k)
frame_vm_group_bin_8127 = frame (4k)
frame_vm_group_bin_8128 = frame (4k)
frame_vm_group_bin_8129 = frame (4k)
frame_vm_group_bin_8130 = frame (4k)
frame_vm_group_bin_8131 = frame (4k)
frame_vm_group_bin_8132 = frame (4k)
frame_vm_group_bin_8133 = frame (4k)
frame_vm_group_bin_8134 = frame (4k)
frame_vm_group_bin_8135 = frame (4k)
frame_vm_group_bin_8136 = frame (4k)
frame_vm_group_bin_8137 = frame (4k)
frame_vm_group_bin_8138 = frame (4k)
frame_vm_group_bin_8139 = frame (4k)
frame_vm_group_bin_8140 = frame (4k)
frame_vm_group_bin_8141 = frame (4k)
frame_vm_group_bin_8142 = frame (4k)
frame_vm_group_bin_8143 = frame (4k)
frame_vm_group_bin_8144 = frame (4k)
frame_vm_group_bin_8145 = frame (4k)
frame_vm_group_bin_8146 = frame (4k)
frame_vm_group_bin_8147 = frame (4k)
frame_vm_group_bin_8148 = frame (4k)
frame_vm_group_bin_8149 = frame (4k)
frame_vm_group_bin_8150 = frame (4k)
frame_vm_group_bin_8151 = frame (4k)
frame_vm_group_bin_8152 = frame (4k)
frame_vm_group_bin_8153 = frame (4k)
frame_vm_group_bin_8154 = frame (4k)
frame_vm_group_bin_8155 = frame (4k)
frame_vm_group_bin_8156 = frame (4k)
frame_vm_group_bin_8157 = frame (4k)
frame_vm_group_bin_8158 = frame (4k)
frame_vm_group_bin_8159 = frame (4k)
frame_vm_group_bin_8160 = frame (4k)
frame_vm_group_bin_8161 = frame (4k)
frame_vm_group_bin_8162 = frame (4k)
frame_vm_group_bin_8163 = frame (4k)
frame_vm_group_bin_8164 = frame (4k)
frame_vm_group_bin_8165 = frame (4k)
frame_vm_group_bin_8166 = frame (4k)
frame_vm_group_bin_8167 = frame (4k)
frame_vm_group_bin_8168 = frame (4k)
frame_vm_group_bin_8169 = frame (4k)
frame_vm_group_bin_8170 = frame (4k)
frame_vm_group_bin_8171 = frame (4k)
frame_vm_group_bin_8172 = frame (4k)
frame_vm_group_bin_8173 = frame (4k)
frame_vm_group_bin_8174 = frame (4k)
frame_vm_group_bin_8175 = frame (4k)
frame_vm_group_bin_8176 = frame (4k)
frame_vm_group_bin_8177 = frame (4k)
frame_vm_group_bin_8178 = frame (4k)
frame_vm_group_bin_8179 = frame (4k)
frame_vm_group_bin_8180 = frame (4k)
frame_vm_group_bin_8181 = frame (4k)
frame_vm_group_bin_8182 = frame (4k)
frame_vm_group_bin_8183 = frame (4k)
frame_vm_group_bin_8184 = frame (4k)
frame_vm_group_bin_8185 = frame (4k)
frame_vm_group_bin_8186 = frame (4k)
frame_vm_group_bin_8187 = frame (4k)
frame_vm_group_bin_8188 = frame (4k)
frame_vm_group_bin_8189 = frame (4k)
frame_vm_group_bin_8190 = frame (4k)
frame_vm_group_bin_8191 = frame (4k)
frame_vm_group_bin_8192 = frame (4k)
frame_vm_group_bin_8193 = frame (4k)
frame_vm_group_bin_8194 = frame (4k)
frame_vm_group_bin_8195 = frame (4k)
frame_vm_group_bin_8196 = frame (4k)
frame_vm_group_bin_8197 = frame (4k)
frame_vm_group_bin_8198 = frame (4k)
frame_vm_group_bin_8199 = frame (4k)
frame_vm_group_bin_8200 = frame (4k)
frame_vm_group_bin_8201 = frame (4k)
frame_vm_group_bin_8202 = frame (4k)
frame_vm_group_bin_8203 = frame (4k)
frame_vm_group_bin_8204 = frame (4k)
frame_vm_group_bin_8205 = frame (4k)
frame_vm_group_bin_8206 = frame (4k)
frame_vm_group_bin_8207 = frame (4k)
frame_vm_group_bin_8208 = frame (4k)
frame_vm_group_bin_8209 = frame (4k)
frame_vm_group_bin_8210 = frame (4k)
frame_vm_group_bin_8211 = frame (4k)
frame_vm_group_bin_8212 = frame (4k)
frame_vm_group_bin_8213 = frame (4k)
frame_vm_group_bin_8214 = frame (4k)
frame_vm_group_bin_8215 = frame (4k)
frame_vm_group_bin_8216 = frame (4k)
frame_vm_group_bin_8217 = frame (4k)
frame_vm_group_bin_8218 = frame (4k)
frame_vm_group_bin_8219 = frame (4k)
frame_vm_group_bin_8220 = frame (4k)
frame_vm_group_bin_8221 = frame (4k)
frame_vm_group_bin_8222 = frame (4k)
frame_vm_group_bin_8223 = frame (4k)
frame_vm_group_bin_8224 = frame (4k)
frame_vm_group_bin_8225 = frame (4k)
frame_vm_group_bin_8226 = frame (4k)
frame_vm_group_bin_8227 = frame (4k)
frame_vm_group_bin_8228 = frame (4k)
frame_vm_group_bin_8229 = frame (4k)
frame_vm_group_bin_8230 = frame (4k)
frame_vm_group_bin_8231 = frame (4k)
frame_vm_group_bin_8232 = frame (4k)
frame_vm_group_bin_8233 = frame (4k)
frame_vm_group_bin_8234 = frame (4k)
frame_vm_group_bin_8235 = frame (4k)
frame_vm_group_bin_8236 = frame (4k)
frame_vm_group_bin_8237 = frame (4k)
frame_vm_group_bin_8238 = frame (4k)
frame_vm_group_bin_8239 = frame (4k)
frame_vm_group_bin_8240 = frame (4k)
frame_vm_group_bin_8241 = frame (4k)
frame_vm_group_bin_8242 = frame (4k)
frame_vm_group_bin_8243 = frame (4k)
frame_vm_group_bin_8244 = frame (4k)
frame_vm_group_bin_8245 = frame (4k)
frame_vm_group_bin_8246 = frame (4k)
frame_vm_group_bin_8247 = frame (4k)
frame_vm_group_bin_8248 = frame (4k)
frame_vm_group_bin_8249 = frame (4k)
frame_vm_group_bin_8250 = frame (4k)
frame_vm_group_bin_8251 = frame (4k)
frame_vm_group_bin_8252 = frame (4k)
frame_vm_group_bin_8253 = frame (4k)
frame_vm_group_bin_8254 = frame (4k)
frame_vm_group_bin_8255 = frame (4k)
frame_vm_group_bin_8256 = frame (4k)
frame_vm_group_bin_8257 = frame (4k)
frame_vm_group_bin_8258 = frame (4k)
frame_vm_group_bin_8259 = frame (4k)
frame_vm_group_bin_8260 = frame (4k)
frame_vm_group_bin_8261 = frame (4k)
frame_vm_group_bin_8262 = frame (4k)
frame_vm_group_bin_8263 = frame (4k)
frame_vm_group_bin_8264 = frame (4k)
frame_vm_group_bin_8265 = frame (4k)
frame_vm_group_bin_8266 = frame (4k)
frame_vm_group_bin_8267 = frame (4k)
frame_vm_group_bin_8268 = frame (4k)
frame_vm_group_bin_8269 = frame (4k)
frame_vm_group_bin_8270 = frame (4k)
frame_vm_group_bin_8271 = frame (4k)
frame_vm_group_bin_8272 = frame (4k)
frame_vm_group_bin_8273 = frame (4k)
frame_vm_group_bin_8274 = frame (4k)
frame_vm_group_bin_8275 = frame (4k)
frame_vm_group_bin_8276 = frame (4k)
frame_vm_group_bin_8277 = frame (4k)
frame_vm_group_bin_8278 = frame (4k)
frame_vm_group_bin_8279 = frame (4k)
frame_vm_group_bin_8280 = frame (4k)
frame_vm_group_bin_8281 = frame (4k)
frame_vm_group_bin_8282 = frame (4k)
frame_vm_group_bin_8283 = frame (4k)
frame_vm_group_bin_8284 = frame (4k)
frame_vm_group_bin_8285 = frame (4k)
frame_vm_group_bin_8286 = frame (4k)
frame_vm_group_bin_8287 = frame (4k)
frame_vm_group_bin_8288 = frame (4k)
frame_vm_group_bin_8289 = frame (4k)
frame_vm_group_bin_8290 = frame (4k)
frame_vm_group_bin_8291 = frame (4k)
frame_vm_group_bin_8292 = frame (4k)
frame_vm_group_bin_8293 = frame (4k)
frame_vm_group_bin_8294 = frame (4k)
frame_vm_group_bin_8295 = frame (4k)
frame_vm_group_bin_8296 = frame (4k)
frame_vm_group_bin_8297 = frame (4k)
frame_vm_group_bin_8298 = frame (4k)
frame_vm_group_bin_8299 = frame (4k)
frame_vm_group_bin_8300 = frame (4k)
frame_vm_group_bin_8301 = frame (4k)
frame_vm_group_bin_8302 = frame (4k)
frame_vm_group_bin_8303 = frame (4k)
frame_vm_group_bin_8304 = frame (4k)
frame_vm_group_bin_8305 = frame (4k)
frame_vm_group_bin_8306 = frame (4k)
frame_vm_group_bin_8307 = frame (4k)
frame_vm_group_bin_8308 = frame (4k)
frame_vm_group_bin_8309 = frame (4k)
frame_vm_group_bin_8310 = frame (4k)
frame_vm_group_bin_8311 = frame (4k)
frame_vm_group_bin_8312 = frame (4k)
frame_vm_group_bin_8313 = frame (4k)
frame_vm_group_bin_8314 = frame (4k)
frame_vm_group_bin_8315 = frame (4k)
frame_vm_group_bin_8316 = frame (4k)
frame_vm_group_bin_8317 = frame (4k)
frame_vm_group_bin_8318 = frame (4k)
frame_vm_group_bin_8319 = frame (4k)
frame_vm_group_bin_8320 = frame (4k)
frame_vm_group_bin_8321 = frame (4k)
frame_vm_group_bin_8322 = frame (4k)
frame_vm_group_bin_8323 = frame (4k)
frame_vm_group_bin_8324 = frame (4k)
frame_vm_group_bin_8325 = frame (4k)
frame_vm_group_bin_8326 = frame (4k)
frame_vm_group_bin_8327 = frame (4k)
frame_vm_group_bin_8328 = frame (4k)
frame_vm_group_bin_8329 = frame (4k)
frame_vm_group_bin_8330 = frame (4k)
frame_vm_group_bin_8331 = frame (4k)
frame_vm_group_bin_8332 = frame (4k)
frame_vm_group_bin_8333 = frame (4k)
frame_vm_group_bin_8334 = frame (4k)
frame_vm_group_bin_8335 = frame (4k)
frame_vm_group_bin_8336 = frame (4k)
frame_vm_group_bin_8337 = frame (4k)
frame_vm_group_bin_8338 = frame (4k)
frame_vm_group_bin_8339 = frame (4k)
frame_vm_group_bin_8340 = frame (4k)
frame_vm_group_bin_8341 = frame (4k)
frame_vm_group_bin_8342 = frame (4k)
frame_vm_group_bin_8343 = frame (4k)
frame_vm_group_bin_8344 = frame (4k)
frame_vm_group_bin_8345 = frame (4k)
frame_vm_group_bin_8346 = frame (4k)
frame_vm_group_bin_8347 = frame (4k)
frame_vm_group_bin_8348 = frame (4k)
frame_vm_group_bin_8349 = frame (4k)
frame_vm_group_bin_8350 = frame (4k)
frame_vm_group_bin_8351 = frame (4k)
frame_vm_group_bin_8352 = frame (4k)
frame_vm_group_bin_8353 = frame (4k)
frame_vm_group_bin_8354 = frame (4k)
frame_vm_group_bin_8355 = frame (4k)
frame_vm_group_bin_8356 = frame (4k)
frame_vm_group_bin_8357 = frame (4k)
frame_vm_group_bin_8358 = frame (4k)
frame_vm_group_bin_8359 = frame (4k)
frame_vm_group_bin_8360 = frame (4k)
frame_vm_group_bin_8361 = frame (4k)
frame_vm_group_bin_8362 = frame (4k)
frame_vm_group_bin_8363 = frame (4k)
frame_vm_group_bin_8364 = frame (4k)
frame_vm_group_bin_8365 = frame (4k)
frame_vm_group_bin_8366 = frame (4k)
frame_vm_group_bin_8367 = frame (4k)
frame_vm_group_bin_8368 = frame (4k)
frame_vm_group_bin_8369 = frame (4k)
frame_vm_group_bin_8370 = frame (4k)
frame_vm_group_bin_8371 = frame (4k)
frame_vm_group_bin_8372 = frame (4k)
frame_vm_group_bin_8373 = frame (4k)
frame_vm_group_bin_8374 = frame (4k)
frame_vm_group_bin_8375 = frame (4k)
frame_vm_group_bin_8376 = frame (4k)
frame_vm_group_bin_8377 = frame (4k)
frame_vm_group_bin_8378 = frame (4k)
frame_vm_group_bin_8379 = frame (4k)
frame_vm_group_bin_8380 = frame (4k)
frame_vm_group_bin_8381 = frame (4k)
frame_vm_group_bin_8382 = frame (4k)
frame_vm_group_bin_8383 = frame (4k)
frame_vm_group_bin_8384 = frame (4k)
frame_vm_group_bin_8385 = frame (4k)
frame_vm_group_bin_8386 = frame (4k)
frame_vm_group_bin_8387 = frame (4k)
frame_vm_group_bin_8388 = frame (4k)
frame_vm_group_bin_8389 = frame (4k)
frame_vm_group_bin_8390 = frame (4k)
frame_vm_group_bin_8391 = frame (4k)
frame_vm_group_bin_8392 = frame (4k)
frame_vm_group_bin_8393 = frame (4k)
frame_vm_group_bin_8394 = frame (4k)
frame_vm_group_bin_8395 = frame (4k)
frame_vm_group_bin_8396 = frame (4k)
frame_vm_group_bin_8397 = frame (4k)
frame_vm_group_bin_8398 = frame (4k)
frame_vm_group_bin_8399 = frame (4k)
frame_vm_group_bin_8400 = frame (4k)
frame_vm_group_bin_8401 = frame (4k)
frame_vm_group_bin_8402 = frame (4k)
frame_vm_group_bin_8403 = frame (4k)
frame_vm_group_bin_8404 = frame (4k)
frame_vm_group_bin_8405 = frame (4k)
frame_vm_group_bin_8406 = frame (4k)
frame_vm_group_bin_8407 = frame (4k)
frame_vm_group_bin_8408 = frame (4k)
frame_vm_group_bin_8409 = frame (4k)
frame_vm_group_bin_8410 = frame (4k)
frame_vm_group_bin_8411 = frame (4k)
frame_vm_group_bin_8412 = frame (4k)
frame_vm_group_bin_8413 = frame (4k)
frame_vm_group_bin_8414 = frame (4k)
frame_vm_group_bin_8415 = frame (4k)
frame_vm_group_bin_8416 = frame (4k)
frame_vm_group_bin_8417 = frame (4k)
frame_vm_group_bin_8418 = frame (4k)
frame_vm_group_bin_8419 = frame (4k)
frame_vm_group_bin_8420 = frame (4k)
frame_vm_group_bin_8421 = frame (4k)
frame_vm_group_bin_8422 = frame (4k)
frame_vm_group_bin_8423 = frame (4k)
frame_vm_group_bin_8424 = frame (4k)
frame_vm_group_bin_8425 = frame (4k)
frame_vm_group_bin_8426 = frame (4k)
frame_vm_group_bin_8427 = frame (4k)
frame_vm_group_bin_8428 = frame (4k)
frame_vm_group_bin_8429 = frame (4k)
frame_vm_group_bin_8430 = frame (4k)
frame_vm_group_bin_8431 = frame (4k)
frame_vm_group_bin_8432 = frame (4k)
frame_vm_group_bin_8433 = frame (4k)
frame_vm_group_bin_8434 = frame (4k)
frame_vm_group_bin_8435 = frame (4k)
frame_vm_group_bin_8436 = frame (4k)
frame_vm_group_bin_8437 = frame (4k)
frame_vm_group_bin_8438 = frame (4k)
frame_vm_group_bin_8439 = frame (4k)
frame_vm_group_bin_8440 = frame (4k)
frame_vm_group_bin_8441 = frame (4k)
frame_vm_group_bin_8442 = frame (4k)
frame_vm_group_bin_8443 = frame (4k)
frame_vm_group_bin_8444 = frame (4k)
frame_vm_group_bin_8445 = frame (4k)
frame_vm_group_bin_8446 = frame (4k)
frame_vm_group_bin_8447 = frame (4k)
frame_vm_group_bin_8448 = frame (4k)
frame_vm_group_bin_8449 = frame (4k)
frame_vm_group_bin_8450 = frame (4k)
frame_vm_group_bin_8451 = frame (4k)
frame_vm_group_bin_8452 = frame (4k)
frame_vm_group_bin_8453 = frame (4k)
frame_vm_group_bin_8454 = frame (4k)
frame_vm_group_bin_8455 = frame (4k)
frame_vm_group_bin_8456 = frame (4k)
frame_vm_group_bin_8457 = frame (4k)
frame_vm_group_bin_8458 = frame (4k)
frame_vm_group_bin_8459 = frame (4k)
frame_vm_group_bin_8460 = frame (4k)
frame_vm_group_bin_8461 = frame (4k)
frame_vm_group_bin_8462 = frame (4k)
frame_vm_group_bin_8463 = frame (4k)
frame_vm_group_bin_8464 = frame (4k)
frame_vm_group_bin_8465 = frame (4k)
frame_vm_group_bin_8466 = frame (4k)
frame_vm_group_bin_8467 = frame (4k)
frame_vm_group_bin_8468 = frame (4k)
frame_vm_group_bin_8469 = frame (4k)
frame_vm_group_bin_8470 = frame (4k)
frame_vm_group_bin_8471 = frame (4k)
frame_vm_group_bin_8472 = frame (4k)
frame_vm_group_bin_8473 = frame (4k)
frame_vm_group_bin_8474 = frame (4k)
frame_vm_group_bin_8475 = frame (4k)
frame_vm_group_bin_8476 = frame (4k)
frame_vm_group_bin_8477 = frame (4k)
frame_vm_group_bin_8478 = frame (4k)
frame_vm_group_bin_8479 = frame (4k)
frame_vm_group_bin_8480 = frame (4k)
frame_vm_group_bin_8481 = frame (4k)
frame_vm_group_bin_8482 = frame (4k)
frame_vm_group_bin_8483 = frame (4k)
frame_vm_group_bin_8484 = frame (4k)
frame_vm_group_bin_8485 = frame (4k)
frame_vm_group_bin_8486 = frame (4k)
frame_vm_group_bin_8487 = frame (4k)
frame_vm_group_bin_8488 = frame (4k)
frame_vm_group_bin_8489 = frame (4k)
frame_vm_group_bin_8490 = frame (4k)
frame_vm_group_bin_8491 = frame (4k)
frame_vm_group_bin_8492 = frame (4k)
frame_vm_group_bin_8493 = frame (4k)
frame_vm_group_bin_8494 = frame (4k)
frame_vm_group_bin_8495 = frame (4k)
frame_vm_group_bin_8496 = frame (4k)
frame_vm_group_bin_8497 = frame (4k)
frame_vm_group_bin_8498 = frame (4k)
frame_vm_group_bin_8499 = frame (4k)
frame_vm_group_bin_8500 = frame (4k)
frame_vm_group_bin_8501 = frame (4k)
frame_vm_group_bin_8502 = frame (4k)
frame_vm_group_bin_8503 = frame (4k)
frame_vm_group_bin_8504 = frame (4k)
frame_vm_group_bin_8505 = frame (4k)
frame_vm_group_bin_8506 = frame (4k)
frame_vm_group_bin_8507 = frame (4k)
frame_vm_group_bin_8508 = frame (4k)
frame_vm_group_bin_8509 = frame (4k)
frame_vm_group_bin_8510 = frame (4k)
frame_vm_group_bin_8511 = frame (4k)
frame_vm_group_bin_8512 = frame (4k)
frame_vm_group_bin_8513 = frame (4k)
frame_vm_group_bin_8514 = frame (4k)
frame_vm_group_bin_8515 = frame (4k)
frame_vm_group_bin_8516 = frame (4k)
frame_vm_group_bin_8517 = frame (4k)
frame_vm_group_bin_8518 = frame (4k)
frame_vm_group_bin_8519 = frame (4k)
frame_vm_group_bin_8520 = frame (4k)
frame_vm_group_bin_8521 = frame (4k)
frame_vm_group_bin_8522 = frame (4k)
frame_vm_group_bin_8523 = frame (4k)
frame_vm_group_bin_8524 = frame (4k)
frame_vm_group_bin_8525 = frame (4k)
frame_vm_group_bin_8526 = frame (4k)
frame_vm_group_bin_8527 = frame (4k)
frame_vm_group_bin_8528 = frame (4k)
frame_vm_group_bin_8529 = frame (4k)
frame_vm_group_bin_8530 = frame (4k)
frame_vm_group_bin_8531 = frame (4k)
frame_vm_group_bin_8532 = frame (4k)
frame_vm_group_bin_8533 = frame (4k)
frame_vm_group_bin_8534 = frame (4k)
frame_vm_group_bin_8535 = frame (4k)
frame_vm_group_bin_8536 = frame (4k)
frame_vm_group_bin_8537 = frame (4k)
frame_vm_group_bin_8538 = frame (4k)
frame_vm_group_bin_8539 = frame (4k)
frame_vm_group_bin_8540 = frame (4k)
frame_vm_group_bin_8541 = frame (4k)
frame_vm_group_bin_8542 = frame (4k)
frame_vm_group_bin_8543 = frame (4k)
frame_vm_group_bin_8544 = frame (4k)
frame_vm_group_bin_8545 = frame (4k)
frame_vm_group_bin_8546 = frame (4k)
frame_vm_group_bin_8547 = frame (4k)
frame_vm_group_bin_8548 = frame (4k)
frame_vm_group_bin_8549 = frame (4k)
frame_vm_group_bin_8550 = frame (4k)
frame_vm_group_bin_8551 = frame (4k)
frame_vm_group_bin_8552 = frame (4k)
frame_vm_group_bin_8553 = frame (4k)
frame_vm_group_bin_8554 = frame (4k)
frame_vm_group_bin_8555 = frame (4k)
frame_vm_group_bin_8556 = frame (4k)
frame_vm_group_bin_8557 = frame (4k)
frame_vm_group_bin_8558 = frame (4k)
frame_vm_group_bin_8559 = frame (4k)
frame_vm_group_bin_8560 = frame (4k)
frame_vm_group_bin_8561 = frame (4k)
frame_vm_group_bin_8562 = frame (4k)
frame_vm_group_bin_8563 = frame (4k)
frame_vm_group_bin_8564 = frame (4k)
frame_vm_group_bin_8565 = frame (4k)
frame_vm_group_bin_8566 = frame (4k)
frame_vm_group_bin_8567 = frame (4k)
frame_vm_group_bin_8568 = frame (4k)
frame_vm_group_bin_8569 = frame (4k)
frame_vm_group_bin_8570 = frame (4k)
frame_vm_group_bin_8571 = frame (4k)
frame_vm_group_bin_8572 = frame (4k)
frame_vm_group_bin_8573 = frame (4k)
frame_vm_group_bin_8574 = frame (4k)
frame_vm_group_bin_8575 = frame (4k)
frame_vm_group_bin_8576 = frame (4k)
frame_vm_group_bin_8577 = frame (4k)
frame_vm_group_bin_8578 = frame (4k)
frame_vm_group_bin_8579 = frame (4k)
frame_vm_group_bin_8580 = frame (4k)
frame_vm_group_bin_8581 = frame (4k)
frame_vm_group_bin_8582 = frame (4k)
frame_vm_group_bin_8583 = frame (4k)
frame_vm_group_bin_8584 = frame (4k)
frame_vm_group_bin_8585 = frame (4k)
frame_vm_group_bin_8586 = frame (4k)
frame_vm_group_bin_8587 = frame (4k)
frame_vm_group_bin_8588 = frame (4k)
frame_vm_group_bin_8589 = frame (4k)
frame_vm_group_bin_8590 = frame (4k)
frame_vm_group_bin_8591 = frame (4k)
frame_vm_group_bin_8592 = frame (4k)
frame_vm_group_bin_8593 = frame (4k)
frame_vm_group_bin_8594 = frame (4k)
frame_vm_group_bin_8595 = frame (4k)
frame_vm_group_bin_8596 = frame (4k)
frame_vm_group_bin_8597 = frame (4k)
frame_vm_group_bin_8598 = frame (4k)
frame_vm_group_bin_8599 = frame (4k)
frame_vm_group_bin_8600 = frame (4k)
frame_vm_group_bin_8601 = frame (4k)
frame_vm_group_bin_8602 = frame (4k)
frame_vm_group_bin_8603 = frame (4k)
frame_vm_group_bin_8604 = frame (4k)
frame_vm_group_bin_8605 = frame (4k)
frame_vm_group_bin_8606 = frame (4k)
frame_vm_group_bin_8607 = frame (4k)
frame_vm_group_bin_8608 = frame (4k)
frame_vm_group_bin_8609 = frame (4k)
frame_vm_group_bin_8610 = frame (4k)
frame_vm_group_bin_8611 = frame (4k)
frame_vm_group_bin_8612 = frame (4k)
frame_vm_group_bin_8613 = frame (4k)
frame_vm_group_bin_8614 = frame (4k)
frame_vm_group_bin_8615 = frame (4k)
frame_vm_group_bin_8616 = frame (4k)
frame_vm_group_bin_8617 = frame (4k)
frame_vm_group_bin_8618 = frame (4k)
frame_vm_group_bin_8619 = frame (4k)
frame_vm_group_bin_8620 = frame (4k)
frame_vm_group_bin_8621 = frame (4k)
frame_vm_group_bin_8622 = frame (4k)
frame_vm_group_bin_8623 = frame (4k)
frame_vm_group_bin_8624 = frame (4k)
frame_vm_group_bin_8625 = frame (4k)
frame_vm_group_bin_8626 = frame (4k)
frame_vm_group_bin_8627 = frame (4k)
frame_vm_group_bin_8628 = frame (4k)
frame_vm_group_bin_8629 = frame (4k)
frame_vm_group_bin_8630 = frame (4k)
frame_vm_group_bin_8631 = frame (4k)
frame_vm_group_bin_8632 = frame (4k)
frame_vm_group_bin_8633 = frame (4k)
frame_vm_group_bin_8634 = frame (4k)
frame_vm_group_bin_8635 = frame (4k)
frame_vm_group_bin_8636 = frame (4k)
frame_vm_group_bin_8637 = frame (4k)
frame_vm_group_bin_8638 = frame (4k)
frame_vm_group_bin_8639 = frame (4k)
frame_vm_group_bin_8640 = frame (4k)
frame_vm_group_bin_8641 = frame (4k)
frame_vm_group_bin_8642 = frame (4k)
frame_vm_group_bin_8643 = frame (4k)
frame_vm_group_bin_8644 = frame (4k)
frame_vm_group_bin_8645 = frame (4k)
frame_vm_group_bin_8646 = frame (4k)
frame_vm_group_bin_8647 = frame (4k)
frame_vm_group_bin_8648 = frame (4k)
frame_vm_group_bin_8649 = frame (4k)
frame_vm_group_bin_8650 = frame (4k)
frame_vm_group_bin_8651 = frame (4k)
frame_vm_group_bin_8652 = frame (4k)
frame_vm_group_bin_8653 = frame (4k)
frame_vm_group_bin_8654 = frame (4k)
frame_vm_group_bin_8655 = frame (4k)
frame_vm_group_bin_8656 = frame (4k)
frame_vm_group_bin_8657 = frame (4k)
frame_vm_group_bin_8658 = frame (4k)
frame_vm_group_bin_8659 = frame (4k)
frame_vm_group_bin_8660 = frame (4k)
frame_vm_group_bin_8661 = frame (4k)
frame_vm_group_bin_8662 = frame (4k)
frame_vm_group_bin_8663 = frame (4k)
frame_vm_group_bin_8664 = frame (4k)
frame_vm_group_bin_8665 = frame (4k)
frame_vm_group_bin_8666 = frame (4k)
frame_vm_group_bin_8667 = frame (4k)
frame_vm_group_bin_8668 = frame (4k)
frame_vm_group_bin_8669 = frame (4k)
frame_vm_group_bin_8670 = frame (4k)
frame_vm_group_bin_8671 = frame (4k)
frame_vm_group_bin_8672 = frame (4k)
frame_vm_group_bin_8673 = frame (4k)
frame_vm_group_bin_8674 = frame (4k)
frame_vm_group_bin_8675 = frame (4k)
frame_vm_group_bin_8676 = frame (4k)
frame_vm_group_bin_8677 = frame (4k)
frame_vm_group_bin_8678 = frame (4k)
frame_vm_group_bin_8679 = frame (4k)
frame_vm_group_bin_8680 = frame (4k)
frame_vm_group_bin_8681 = frame (4k)
frame_vm_group_bin_8682 = frame (4k)
frame_vm_group_bin_8683 = frame (4k)
frame_vm_group_bin_8684 = frame (4k)
frame_vm_group_bin_8685 = frame (4k)
frame_vm_group_bin_8686 = frame (4k)
frame_vm_group_bin_8687 = frame (4k)
frame_vm_group_bin_8688 = frame (4k)
frame_vm_group_bin_8689 = frame (4k)
frame_vm_group_bin_8690 = frame (4k)
frame_vm_group_bin_8691 = frame (4k)
frame_vm_group_bin_8692 = frame (4k)
frame_vm_group_bin_8693 = frame (4k)
frame_vm_group_bin_8694 = frame (4k)
frame_vm_group_bin_8695 = frame (4k)
frame_vm_group_bin_8696 = frame (4k)
frame_vm_group_bin_8697 = frame (4k)
frame_vm_group_bin_8698 = frame (4k)
frame_vm_group_bin_8699 = frame (4k)
frame_vm_group_bin_8700 = frame (4k)
frame_vm_group_bin_8701 = frame (4k)
frame_vm_group_bin_8702 = frame (4k)
frame_vm_group_bin_8703 = frame (4k)
frame_vm_group_bin_8704 = frame (4k)
frame_vm_group_bin_8705 = frame (4k)
frame_vm_group_bin_8706 = frame (4k)
frame_vm_group_bin_8707 = frame (4k)
frame_vm_group_bin_8708 = frame (4k)
frame_vm_group_bin_8709 = frame (4k)
frame_vm_group_bin_8710 = frame (4k)
frame_vm_group_bin_8711 = frame (4k)
frame_vm_group_bin_8712 = frame (4k)
frame_vm_group_bin_8713 = frame (4k)
frame_vm_group_bin_8714 = frame (4k)
frame_vm_group_bin_8715 = frame (4k)
frame_vm_group_bin_8716 = frame (4k)
frame_vm_group_bin_8717 = frame (4k)
frame_vm_group_bin_8718 = frame (4k)
frame_vm_group_bin_8719 = frame (4k)
frame_vm_group_bin_8720 = frame (4k)
frame_vm_group_bin_8721 = frame (4k)
frame_vm_group_bin_8722 = frame (4k)
frame_vm_group_bin_8723 = frame (4k)
frame_vm_group_bin_8724 = frame (4k)
frame_vm_group_bin_8725 = frame (4k)
frame_vm_group_bin_8726 = frame (4k)
frame_vm_group_bin_8727 = frame (4k)
frame_vm_group_bin_8728 = frame (4k)
frame_vm_group_bin_8729 = frame (4k)
frame_vm_group_bin_8730 = frame (4k)
frame_vm_group_bin_8731 = frame (4k)
frame_vm_group_bin_8732 = frame (4k)
frame_vm_group_bin_8733 = frame (4k)
frame_vm_group_bin_8734 = frame (4k)
frame_vm_group_bin_8735 = frame (4k)
frame_vm_group_bin_8736 = frame (4k)
frame_vm_group_bin_8737 = frame (4k)
frame_vm_group_bin_8738 = frame (4k)
frame_vm_group_bin_8739 = frame (4k)
frame_vm_group_bin_8740 = frame (4k)
frame_vm_group_bin_8741 = frame (4k)
frame_vm_group_bin_8742 = frame (4k)
frame_vm_group_bin_8743 = frame (4k)
frame_vm_group_bin_8744 = frame (4k)
frame_vm_group_bin_8745 = frame (4k)
frame_vm_group_bin_8746 = frame (4k)
frame_vm_group_bin_8747 = frame (4k)
frame_vm_group_bin_8748 = frame (4k)
frame_vm_group_bin_8749 = frame (4k)
frame_vm_group_bin_8750 = frame (4k)
frame_vm_group_bin_8751 = frame (4k)
frame_vm_group_bin_8752 = frame (4k)
frame_vm_group_bin_8753 = frame (4k)
frame_vm_group_bin_8754 = frame (4k)
frame_vm_group_bin_8755 = frame (4k)
frame_vm_group_bin_8756 = frame (4k)
frame_vm_group_bin_8757 = frame (4k)
frame_vm_group_bin_8758 = frame (4k)
frame_vm_group_bin_8759 = frame (4k)
frame_vm_group_bin_8760 = frame (4k)
frame_vm_group_bin_8761 = frame (4k)
frame_vm_group_bin_8762 = frame (4k)
frame_vm_group_bin_8763 = frame (4k)
frame_vm_group_bin_8764 = frame (4k)
frame_vm_group_bin_8765 = frame (4k)
frame_vm_group_bin_8766 = frame (4k)
frame_vm_group_bin_8767 = frame (4k)
frame_vm_group_bin_8768 = frame (4k)
frame_vm_group_bin_8769 = frame (4k)
frame_vm_group_bin_8770 = frame (4k)
frame_vm_group_bin_8771 = frame (4k)
frame_vm_group_bin_8772 = frame (4k)
frame_vm_group_bin_8773 = frame (4k)
frame_vm_group_bin_8774 = frame (4k)
frame_vm_group_bin_8775 = frame (4k)
frame_vm_group_bin_8776 = frame (4k)
frame_vm_group_bin_8777 = frame (4k)
frame_vm_group_bin_8778 = frame (4k)
frame_vm_group_bin_8779 = frame (4k)
frame_vm_group_bin_8780 = frame (4k)
frame_vm_group_bin_8781 = frame (4k)
frame_vm_group_bin_8782 = frame (4k)
frame_vm_group_bin_8783 = frame (4k)
frame_vm_group_bin_8784 = frame (4k)
frame_vm_group_bin_8785 = frame (4k)
frame_vm_group_bin_8786 = frame (4k)
frame_vm_group_bin_8787 = frame (4k)
frame_vm_group_bin_8788 = frame (4k)
frame_vm_group_bin_8789 = frame (4k)
frame_vm_group_bin_8790 = frame (4k)
frame_vm_group_bin_8791 = frame (4k)
frame_vm_group_bin_8792 = frame (4k)
frame_vm_group_bin_8793 = frame (4k)
frame_vm_group_bin_8794 = frame (4k)
frame_vm_group_bin_8795 = frame (4k)
frame_vm_group_bin_8796 = frame (4k)
frame_vm_group_bin_8797 = frame (4k)
frame_vm_group_bin_8798 = frame (4k)
frame_vm_group_bin_8799 = frame (4k)
frame_vm_group_bin_8800 = frame (4k)
frame_vm_group_bin_8801 = frame (4k)
frame_vm_group_bin_8802 = frame (4k)
frame_vm_group_bin_8803 = frame (4k)
frame_vm_group_bin_8804 = frame (4k)
frame_vm_group_bin_8805 = frame (4k)
frame_vm_group_bin_8806 = frame (4k)
frame_vm_group_bin_8807 = frame (4k)
frame_vm_group_bin_8808 = frame (4k)
frame_vm_group_bin_8809 = frame (4k)
frame_vm_group_bin_8810 = frame (4k)
frame_vm_group_bin_8811 = frame (4k)
frame_vm_group_bin_8812 = frame (4k)
frame_vm_group_bin_8813 = frame (4k)
frame_vm_group_bin_8814 = frame (4k)
frame_vm_group_bin_8815 = frame (4k)
frame_vm_group_bin_8816 = frame (4k)
frame_vm_group_bin_8817 = frame (4k)
frame_vm_group_bin_8818 = frame (4k)
frame_vm_group_bin_8819 = frame (4k)
frame_vm_group_bin_8820 = frame (4k)
frame_vm_group_bin_8821 = frame (4k)
frame_vm_group_bin_8822 = frame (4k)
frame_vm_group_bin_8823 = frame (4k)
frame_vm_group_bin_8824 = frame (4k)
frame_vm_group_bin_8825 = frame (4k)
frame_vm_group_bin_8826 = frame (4k)
frame_vm_group_bin_8827 = frame (4k)
frame_vm_group_bin_8828 = frame (4k)
frame_vm_group_bin_8829 = frame (4k)
frame_vm_group_bin_8830 = frame (4k)
frame_vm_group_bin_8831 = frame (4k)
frame_vm_group_bin_8832 = frame (4k)
frame_vm_group_bin_8833 = frame (4k)
frame_vm_group_bin_8834 = frame (4k)
frame_vm_group_bin_8835 = frame (4k)
frame_vm_group_bin_8836 = frame (4k)
frame_vm_group_bin_8837 = frame (4k)
frame_vm_group_bin_8838 = frame (4k)
frame_vm_group_bin_8839 = frame (4k)
frame_vm_group_bin_8840 = frame (4k)
frame_vm_group_bin_8841 = frame (4k)
frame_vm_group_bin_8842 = frame (4k)
frame_vm_group_bin_8843 = frame (4k)
frame_vm_group_bin_8844 = frame (4k)
frame_vm_group_bin_8845 = frame (4k)
frame_vm_group_bin_8846 = frame (4k)
frame_vm_group_bin_8847 = frame (4k)
frame_vm_group_bin_8848 = frame (4k)
frame_vm_group_bin_8849 = frame (4k)
frame_vm_group_bin_8850 = frame (4k)
frame_vm_group_bin_8851 = frame (4k)
frame_vm_group_bin_8852 = frame (4k)
frame_vm_group_bin_8853 = frame (4k)
frame_vm_group_bin_8854 = frame (4k)
frame_vm_group_bin_8856 = frame (4k)
frame_vm_group_bin_8857 = frame (4k)
frame_vm_group_bin_8858 = frame (4k)
frame_vm_group_bin_8859 = frame (4k)
frame_vm_group_bin_8860 = frame (4k)
frame_vm_group_bin_8861 = frame (4k)
frame_vm_group_bin_8862 = frame (4k)
frame_vm_group_bin_8863 = frame (4k)
frame_vm_group_bin_8864 = frame (4k)
frame_vm_group_bin_8865 = frame (4k)
frame_vm_group_bin_8866 = frame (4k)
frame_vm_group_bin_8867 = frame (4k)
frame_vm_group_bin_8868 = frame (4k)
frame_vm_group_bin_8869 = frame (4k)
frame_vm_group_bin_8870 = frame (4k)
frame_vm_group_bin_8871 = frame (4k)
frame_vm_group_bin_8872 = frame (4k)
frame_vm_group_bin_8873 = frame (4k)
frame_vm_group_bin_8874 = frame (4k)
frame_vm_group_bin_8875 = frame (4k)
frame_vm_group_bin_8876 = frame (4k)
frame_vm_group_bin_8877 = frame (4k)
frame_vm_group_bin_8878 = frame (4k)
frame_vm_group_bin_8879 = frame (4k)
frame_vm_group_bin_8880 = frame (4k)
frame_vm_group_bin_8881 = frame (4k)
frame_vm_group_bin_8882 = frame (4k)
frame_vm_group_bin_8883 = frame (4k)
frame_vm_group_bin_8884 = frame (4k)
frame_vm_group_bin_8885 = frame (4k)
frame_vm_group_bin_8886 = frame (4k)
frame_vm_group_bin_8887 = frame (4k)
frame_vm_group_bin_8888 = frame (4k)
frame_vm_group_bin_8889 = frame (4k)
frame_vm_group_bin_8890 = frame (4k)
frame_vm_group_bin_8891 = frame (4k)
frame_vm_group_bin_8892 = frame (4k)
frame_vm_group_bin_8893 = frame (4k)
frame_vm_group_bin_8894 = frame (4k)
frame_vm_group_bin_8895 = frame (4k)
frame_vm_group_bin_8896 = frame (4k)
frame_vm_group_bin_8897 = frame (4k)
frame_vm_group_bin_8898 = frame (4k)
frame_vm_group_bin_8899 = frame (4k)
frame_vm_group_bin_8900 = frame (4k)
frame_vm_group_bin_8901 = frame (4k)
frame_vm_group_bin_8902 = frame (4k)
frame_vm_group_bin_8903 = frame (4k)
frame_vm_group_bin_8904 = frame (4k)
frame_vm_group_bin_8905 = frame (4k)
frame_vm_group_bin_8906 = frame (4k)
frame_vm_group_bin_8907 = frame (4k)
frame_vm_group_bin_8908 = frame (4k)
frame_vm_group_bin_8909 = frame (4k)
frame_vm_group_bin_8910 = frame (4k)
frame_vm_group_bin_8911 = frame (4k)
frame_vm_group_bin_8912 = frame (4k)
frame_vm_group_bin_8913 = frame (4k)
frame_vm_group_bin_8914 = frame (4k)
frame_vm_group_bin_8915 = frame (4k)
frame_vm_group_bin_8916 = frame (4k)
frame_vm_group_bin_8917 = frame (4k)
frame_vm_group_bin_8918 = frame (4k)
frame_vm_group_bin_8919 = frame (4k)
frame_vm_group_bin_8920 = frame (4k)
frame_vm_group_bin_8921 = frame (4k)
frame_vm_group_bin_8922 = frame (4k)
frame_vm_group_bin_8923 = frame (4k)
frame_vm_group_bin_8924 = frame (4k)
frame_vm_group_bin_8925 = frame (4k)
frame_vm_group_bin_8926 = frame (4k)
frame_vm_group_bin_8927 = frame (4k)
frame_vm_group_bin_8928 = frame (4k)
frame_vm_group_bin_8929 = frame (4k)
frame_vm_group_bin_8930 = frame (4k)
frame_vm_group_bin_8931 = frame (4k)
frame_vm_group_bin_8932 = frame (4k)
frame_vm_group_bin_8933 = frame (4k)
frame_vm_group_bin_8934 = frame (4k)
frame_vm_group_bin_8935 = frame (4k)
frame_vm_group_bin_8936 = frame (4k)
frame_vm_group_bin_8937 = frame (4k)
frame_vm_group_bin_8938 = frame (4k)
frame_vm_group_bin_8939 = frame (4k)
frame_vm_group_bin_8940 = frame (4k)
frame_vm_group_bin_8941 = frame (4k)
frame_vm_group_bin_8942 = frame (4k)
frame_vm_group_bin_8943 = frame (4k)
frame_vm_group_bin_8944 = frame (4k)
frame_vm_group_bin_8945 = frame (4k)
frame_vm_group_bin_8946 = frame (4k)
frame_vm_group_bin_8947 = frame (4k)
frame_vm_group_bin_8948 = frame (4k)
frame_vm_group_bin_8949 = frame (4k)
frame_vm_group_bin_8950 = frame (4k)
frame_vm_group_bin_8951 = frame (4k)
frame_vm_group_bin_8952 = frame (4k)
frame_vm_group_bin_8953 = frame (4k)
frame_vm_group_bin_8954 = frame (4k)
frame_vm_group_bin_8955 = frame (4k)
frame_vm_group_bin_8956 = frame (4k)
frame_vm_group_bin_8957 = frame (4k)
frame_vm_group_bin_8958 = frame (4k)
frame_vm_group_bin_8959 = frame (4k)
frame_vm_group_bin_8960 = frame (4k)
frame_vm_group_bin_8961 = frame (4k)
frame_vm_group_bin_8962 = frame (4k)
frame_vm_group_bin_8963 = frame (4k)
frame_vm_group_bin_8964 = frame (4k)
frame_vm_group_bin_8965 = frame (4k)
frame_vm_group_bin_8966 = frame (4k)
frame_vm_group_bin_8967 = frame (4k)
frame_vm_group_bin_8968 = frame (4k)
frame_vm_group_bin_8969 = frame (4k)
frame_vm_group_bin_8970 = frame (4k)
frame_vm_group_bin_8971 = frame (4k)
frame_vm_group_bin_8972 = frame (4k)
frame_vm_group_bin_8973 = frame (4k)
frame_vm_group_bin_8974 = frame (4k)
frame_vm_group_bin_8975 = frame (4k)
frame_vm_group_bin_8976 = frame (4k)
frame_vm_group_bin_8977 = frame (4k)
frame_vm_group_bin_8978 = frame (4k)
frame_vm_group_bin_8979 = frame (4k)
frame_vm_group_bin_8980 = frame (4k)
frame_vm_group_bin_8981 = frame (4k)
frame_vm_group_bin_8982 = frame (4k)
frame_vm_group_bin_8983 = frame (4k)
frame_vm_group_bin_8984 = frame (4k)
frame_vm_group_bin_8985 = frame (4k)
frame_vm_group_bin_8986 = frame (4k)
frame_vm_group_bin_8987 = frame (4k)
frame_vm_group_bin_8988 = frame (4k)
frame_vm_group_bin_8989 = frame (4k)
frame_vm_group_bin_8990 = frame (4k)
frame_vm_group_bin_8991 = frame (4k)
frame_vm_group_bin_8992 = frame (4k)
frame_vm_group_bin_8993 = frame (4k)
frame_vm_group_bin_8994 = frame (4k)
frame_vm_group_bin_8995 = frame (4k)
frame_vm_group_bin_8996 = frame (4k)
frame_vm_group_bin_8997 = frame (4k)
frame_vm_group_bin_8998 = frame (4k)
frame_vm_group_bin_8999 = frame (4k)
frame_vm_group_bin_9000 = frame (4k)
frame_vm_group_bin_9001 = frame (4k)
frame_vm_group_bin_9002 = frame (4k)
frame_vm_group_bin_9003 = frame (4k)
frame_vm_group_bin_9004 = frame (4k)
frame_vm_group_bin_9005 = frame (4k)
frame_vm_group_bin_9006 = frame (4k)
frame_vm_group_bin_9007 = frame (4k)
frame_vm_group_bin_9008 = frame (4k)
frame_vm_group_bin_9009 = frame (4k)
frame_vm_group_bin_9010 = frame (4k)
frame_vm_group_bin_9011 = frame (4k)
frame_vm_group_bin_9012 = frame (4k)
frame_vm_group_bin_9013 = frame (4k)
frame_vm_group_bin_9014 = frame (4k)
frame_vm_group_bin_9015 = frame (4k)
frame_vm_group_bin_9016 = frame (4k)
frame_vm_group_bin_9017 = frame (4k)
frame_vm_group_bin_9018 = frame (4k)
frame_vm_group_bin_9019 = frame (4k)
frame_vm_group_bin_9020 = frame (4k)
frame_vm_group_bin_9021 = frame (4k)
frame_vm_group_bin_9022 = frame (4k)
frame_vm_group_bin_9023 = frame (4k)
frame_vm_group_bin_9024 = frame (4k)
frame_vm_group_bin_9025 = frame (4k)
frame_vm_group_bin_9026 = frame (4k)
frame_vm_group_bin_9027 = frame (4k)
frame_vm_group_bin_9028 = frame (4k)
frame_vm_group_bin_9029 = frame (4k)
frame_vm_group_bin_9030 = frame (4k)
frame_vm_group_bin_9031 = frame (4k)
frame_vm_group_bin_9032 = frame (4k)
frame_vm_group_bin_9033 = frame (4k)
frame_vm_group_bin_9034 = frame (4k)
frame_vm_group_bin_9035 = frame (4k)
frame_vm_group_bin_9036 = frame (4k)
frame_vm_group_bin_9037 = frame (4k)
frame_vm_group_bin_9038 = frame (4k)
frame_vm_group_bin_9039 = frame (4k)
frame_vm_group_bin_9040 = frame (4k)
frame_vm_group_bin_9041 = frame (4k)
frame_vm_group_bin_9042 = frame (4k)
frame_vm_group_bin_9043 = frame (4k)
frame_vm_group_bin_9044 = frame (4k)
frame_vm_group_bin_9045 = frame (4k)
frame_vm_group_bin_9046 = frame (4k)
frame_vm_group_bin_9047 = frame (4k)
frame_vm_group_bin_9048 = frame (4k)
frame_vm_group_bin_9049 = frame (4k)
frame_vm_group_bin_9050 = frame (4k)
frame_vm_group_bin_9051 = frame (4k)
frame_vm_group_bin_9052 = frame (4k)
frame_vm_group_bin_9053 = frame (4k)
frame_vm_group_bin_9054 = frame (4k)
frame_vm_group_bin_9055 = frame (4k)
frame_vm_group_bin_9056 = frame (4k)
frame_vm_group_bin_9057 = frame (4k)
frame_vm_group_bin_9058 = frame (4k)
frame_vm_group_bin_9059 = frame (4k)
frame_vm_group_bin_9060 = frame (4k)
frame_vm_group_bin_9061 = frame (4k)
frame_vm_group_bin_9062 = frame (4k)
frame_vm_group_bin_9063 = frame (4k)
frame_vm_group_bin_9064 = frame (4k)
frame_vm_group_bin_9065 = frame (4k)
frame_vm_group_bin_9066 = frame (4k)
frame_vm_group_bin_9067 = frame (4k)
frame_vm_group_bin_9068 = frame (4k)
frame_vm_group_bin_9069 = frame (4k)
frame_vm_group_bin_9070 = frame (4k)
frame_vm_group_bin_9071 = frame (4k)
frame_vm_group_bin_9072 = frame (4k)
frame_vm_group_bin_9073 = frame (4k)
frame_vm_group_bin_9074 = frame (4k)
frame_vm_group_bin_9075 = frame (4k)
frame_vm_group_bin_9076 = frame (4k)
frame_vm_group_bin_9077 = frame (4k)
frame_vm_group_bin_9078 = frame (4k)
frame_vm_group_bin_9079 = frame (4k)
frame_vm_group_bin_9080 = frame (4k)
frame_vm_group_bin_9081 = frame (4k)
frame_vm_group_bin_9082 = frame (4k)
frame_vm_group_bin_9083 = frame (4k)
frame_vm_group_bin_9084 = frame (4k)
frame_vm_group_bin_9085 = frame (4k)
frame_vm_group_bin_9086 = frame (4k)
frame_vm_group_bin_9087 = frame (4k)
frame_vm_group_bin_9088 = frame (4k)
frame_vm_group_bin_9089 = frame (4k)
frame_vm_group_bin_9090 = frame (4k)
frame_vm_group_bin_9091 = frame (4k)
frame_vm_group_bin_9092 = frame (4k)
frame_vm_group_bin_9093 = frame (4k)
frame_vm_group_bin_9094 = frame (4k)
frame_vm_group_bin_9095 = frame (4k)
frame_vm_group_bin_9096 = frame (4k)
frame_vm_group_bin_9097 = frame (4k)
frame_vm_group_bin_9098 = frame (4k)
frame_vm_group_bin_9099 = frame (4k)
frame_vm_group_bin_9100 = frame (4k)
frame_vm_group_bin_9101 = frame (4k)
frame_vm_group_bin_9102 = frame (4k)
frame_vm_group_bin_9103 = frame (4k)
frame_vm_group_bin_9104 = frame (4k)
frame_vm_group_bin_9105 = frame (4k)
frame_vm_group_bin_9106 = frame (4k)
frame_vm_group_bin_9107 = frame (4k)
frame_vm_group_bin_9108 = frame (4k)
frame_vm_group_bin_9109 = frame (4k)
frame_vm_group_bin_9110 = frame (4k)
frame_vm_group_bin_9111 = frame (4k)
frame_vm_group_bin_9112 = frame (4k)
frame_vm_group_bin_9113 = frame (4k)
frame_vm_group_bin_9114 = frame (4k)
frame_vm_group_bin_9115 = frame (4k)
frame_vm_group_bin_9116 = frame (4k)
frame_vm_group_bin_9117 = frame (4k)
frame_vm_group_bin_9118 = frame (4k)
frame_vm_group_bin_9119 = frame (4k)
frame_vm_group_bin_9120 = frame (4k)
frame_vm_group_bin_9121 = frame (4k)
frame_vm_group_bin_9122 = frame (4k)
frame_vm_group_bin_9123 = frame (4k)
frame_vm_group_bin_9124 = frame (4k)
frame_vm_group_bin_9125 = frame (4k)
frame_vm_group_bin_9126 = frame (4k)
frame_vm_group_bin_9127 = frame (4k)
frame_vm_group_bin_9128 = frame (4k)
frame_vm_group_bin_9129 = frame (4k)
frame_vm_group_bin_9130 = frame (4k)
frame_vm_group_bin_9131 = frame (4k)
frame_vm_group_bin_9132 = frame (4k)
frame_vm_group_bin_9133 = frame (4k)
frame_vm_group_bin_9134 = frame (4k)
frame_vm_group_bin_9135 = frame (4k)
frame_vm_group_bin_9136 = frame (4k)
frame_vm_group_bin_9137 = frame (4k)
frame_vm_group_bin_9138 = frame (4k)
frame_vm_group_bin_9139 = frame (4k)
frame_vm_group_bin_9140 = frame (4k)
frame_vm_group_bin_9141 = frame (4k)
frame_vm_group_bin_9142 = frame (4k)
frame_vm_group_bin_9143 = frame (4k)
frame_vm_group_bin_9144 = frame (4k)
frame_vm_group_bin_9145 = frame (4k)
frame_vm_group_bin_9146 = frame (4k)
frame_vm_group_bin_9147 = frame (4k)
frame_vm_group_bin_9148 = frame (4k)
frame_vm_group_bin_9149 = frame (4k)
frame_vm_group_bin_9150 = frame (4k)
frame_vm_group_bin_9151 = frame (4k)
frame_vm_group_bin_9152 = frame (4k)
frame_vm_group_bin_9153 = frame (4k)
frame_vm_group_bin_9154 = frame (4k)
frame_vm_group_bin_9155 = frame (4k)
frame_vm_group_bin_9156 = frame (4k)
frame_vm_group_bin_9157 = frame (4k)
frame_vm_group_bin_9158 = frame (4k)
frame_vm_group_bin_9159 = frame (4k)
frame_vm_group_bin_9160 = frame (4k)
frame_vm_group_bin_9161 = frame (4k)
frame_vm_group_bin_9162 = frame (4k)
frame_vm_group_bin_9163 = frame (4k)
frame_vm_group_bin_9164 = frame (4k)
frame_vm_group_bin_9165 = frame (4k)
frame_vm_group_bin_9166 = frame (4k)
frame_vm_group_bin_9167 = frame (4k)
frame_vm_group_bin_9168 = frame (4k)
frame_vm_group_bin_9169 = frame (4k)
frame_vm_group_bin_9170 = frame (4k)
frame_vm_group_bin_9171 = frame (4k)
frame_vm_group_bin_9172 = frame (4k)
frame_vm_group_bin_9173 = frame (4k)
frame_vm_group_bin_9174 = frame (4k)
frame_vm_group_bin_9175 = frame (4k)
frame_vm_group_bin_9176 = frame (4k)
frame_vm_group_bin_9177 = frame (4k)
frame_vm_group_bin_9178 = frame (4k)
frame_vm_group_bin_9179 = frame (4k)
frame_vm_group_bin_9180 = frame (4k)
frame_vm_group_bin_9181 = frame (4k)
frame_vm_group_bin_9182 = frame (4k)
frame_vm_group_bin_9183 = frame (4k)
frame_vm_group_bin_9184 = frame (4k)
frame_vm_group_bin_9185 = frame (4k)
frame_vm_group_bin_9186 = frame (4k)
frame_vm_group_bin_9187 = frame (4k)
frame_vm_group_bin_9188 = frame (4k)
frame_vm_group_bin_9189 = frame (4k)
frame_vm_group_bin_9190 = frame (4k)
frame_vm_group_bin_9191 = frame (4k)
frame_vm_group_bin_9192 = frame (4k)
frame_vm_group_bin_9193 = frame (4k)
frame_vm_group_bin_9194 = frame (4k)
frame_vm_group_bin_9195 = frame (4k)
frame_vm_group_bin_9196 = frame (4k)
frame_vm_group_bin_9197 = frame (4k)
frame_vm_group_bin_9198 = frame (4k)
frame_vm_group_bin_9199 = frame (4k)
frame_vm_group_bin_9200 = frame (4k)
frame_vm_group_bin_9201 = frame (4k)
frame_vm_group_bin_9202 = frame (4k)
frame_vm_group_bin_9203 = frame (4k)
frame_vm_group_bin_9204 = frame (4k)
frame_vm_group_bin_9205 = frame (4k)
frame_vm_group_bin_9206 = frame (4k)
frame_vm_group_bin_9207 = frame (4k)
frame_vm_group_bin_9208 = frame (4k)
frame_vm_group_bin_9209 = frame (4k)
frame_vm_group_bin_9210 = frame (4k)
frame_vm_group_bin_9211 = frame (4k)
frame_vm_group_bin_9212 = frame (4k)
frame_vm_group_bin_9213 = frame (4k)
frame_vm_group_bin_9214 = frame (4k)
frame_vm_group_bin_9215 = frame (4k)
frame_vm_group_bin_9216 = frame (4k)
frame_vm_group_bin_9217 = frame (4k)
frame_vm_group_bin_9218 = frame (4k)
frame_vm_group_bin_9219 = frame (4k)
frame_vm_group_bin_9220 = frame (4k)
frame_vm_group_bin_9221 = frame (4k)
frame_vm_group_bin_9222 = frame (4k)
frame_vm_group_bin_9223 = frame (4k)
frame_vm_group_bin_9224 = frame (4k)
frame_vm_group_bin_9225 = frame (4k)
frame_vm_group_bin_9226 = frame (4k)
frame_vm_group_bin_9227 = frame (4k)
frame_vm_group_bin_9228 = frame (4k)
frame_vm_group_bin_9229 = frame (4k)
frame_vm_group_bin_9230 = frame (4k)
frame_vm_group_bin_9231 = frame (4k)
frame_vm_group_bin_9232 = frame (4k)
frame_vm_group_bin_9233 = frame (4k)
frame_vm_group_bin_9234 = frame (4k)
frame_vm_group_bin_9235 = frame (4k)
frame_vm_group_bin_9236 = frame (4k)
frame_vm_group_bin_9237 = frame (4k)
frame_vm_group_bin_9238 = frame (4k)
frame_vm_group_bin_9239 = frame (4k)
frame_vm_group_bin_9240 = frame (4k)
frame_vm_group_bin_9241 = frame (4k)
frame_vm_group_bin_9242 = frame (4k)
frame_vm_group_bin_9243 = frame (4k)
frame_vm_group_bin_9244 = frame (4k)
frame_vm_group_bin_9245 = frame (4k)
frame_vm_group_bin_9246 = frame (4k)
frame_vm_group_bin_9247 = frame (4k)
frame_vm_group_bin_9248 = frame (4k)
frame_vm_group_bin_9249 = frame (4k)
frame_vm_group_bin_9250 = frame (4k)
frame_vm_group_bin_9251 = frame (4k)
frame_vm_group_bin_9252 = frame (4k)
frame_vm_group_bin_9253 = frame (4k)
frame_vm_group_bin_9254 = frame (4k)
frame_vm_group_bin_9255 = frame (4k)
frame_vm_group_bin_9256 = frame (4k)
frame_vm_group_bin_9257 = frame (4k)
frame_vm_group_bin_9258 = frame (4k)
frame_vm_group_bin_9259 = frame (4k)
frame_vm_group_bin_9260 = frame (4k)
frame_vm_group_bin_9261 = frame (4k)
frame_vm_group_bin_9262 = frame (4k)
frame_vm_group_bin_9263 = frame (4k)
frame_vm_group_bin_9264 = frame (4k)
frame_vm_group_bin_9265 = frame (4k)
frame_vm_group_bin_9266 = frame (4k)
frame_vm_group_bin_9267 = frame (4k)
frame_vm_group_bin_9268 = frame (4k)
frame_vm_group_bin_9269 = frame (4k)
frame_vm_group_bin_9270 = frame (4k)
frame_vm_group_bin_9271 = frame (4k)
frame_vm_group_bin_9272 = frame (4k)
frame_vm_group_bin_9273 = frame (4k)
frame_vm_group_bin_9274 = frame (4k)
frame_vm_group_bin_9275 = frame (4k)
frame_vm_group_bin_9276 = frame (4k)
frame_vm_group_bin_9277 = frame (4k)
frame_vm_group_bin_9278 = frame (4k)
frame_vm_group_bin_9279 = frame (4k)
frame_vm_group_bin_9280 = frame (4k)
frame_vm_group_bin_9281 = frame (4k)
frame_vm_group_bin_9282 = frame (4k)
frame_vm_group_bin_9283 = frame (4k)
frame_vm_group_bin_9284 = frame (4k)
frame_vm_group_bin_9285 = frame (4k)
frame_vm_group_bin_9286 = frame (4k)
frame_vm_group_bin_9287 = frame (4k)
frame_vm_group_bin_9288 = frame (4k)
frame_vm_group_bin_9289 = frame (4k)
frame_vm_group_bin_9290 = frame (4k)
frame_vm_group_bin_9291 = frame (4k)
frame_vm_group_bin_9292 = frame (4k)
frame_vm_group_bin_9293 = frame (4k)
frame_vm_group_bin_9294 = frame (4k)
frame_vm_group_bin_9295 = frame (4k)
frame_vm_group_bin_9296 = frame (4k)
frame_vm_group_bin_9297 = frame (4k)
frame_vm_group_bin_9298 = frame (4k)
frame_vm_group_bin_9299 = frame (4k)
frame_vm_group_bin_9300 = frame (4k)
frame_vm_group_bin_9301 = frame (4k)
frame_vm_group_bin_9302 = frame (4k)
frame_vm_group_bin_9303 = frame (4k)
frame_vm_group_bin_9304 = frame (4k)
frame_vm_group_bin_9305 = frame (4k)
frame_vm_group_bin_9306 = frame (4k)
frame_vm_group_bin_9307 = frame (4k)
frame_vm_group_bin_9308 = frame (4k)
frame_vm_group_bin_9309 = frame (4k)
frame_vm_group_bin_9310 = frame (4k)
frame_vm_group_bin_9311 = frame (4k)
frame_vm_group_bin_9312 = frame (4k)
frame_vm_group_bin_9313 = frame (4k)
frame_vm_group_bin_9314 = frame (4k)
frame_vm_group_bin_9315 = frame (4k)
frame_vm_group_bin_9316 = frame (4k)
frame_vm_group_bin_9317 = frame (4k)
frame_vm_group_bin_9318 = frame (4k)
frame_vm_group_bin_9319 = frame (4k)
frame_vm_group_bin_9320 = frame (4k)
frame_vm_group_bin_9321 = frame (4k)
frame_vm_group_bin_9322 = frame (4k)
frame_vm_group_bin_9323 = frame (4k)
frame_vm_group_bin_9324 = frame (4k)
frame_vm_group_bin_9325 = frame (4k)
frame_vm_group_bin_9326 = frame (4k)
frame_vm_group_bin_9327 = frame (4k)
frame_vm_group_bin_9328 = frame (4k)
frame_vm_group_bin_9329 = frame (4k)
frame_vm_group_bin_9330 = frame (4k)
frame_vm_group_bin_9331 = frame (4k)
frame_vm_group_bin_9332 = frame (4k)
frame_vm_group_bin_9333 = frame (4k)
frame_vm_group_bin_9334 = frame (4k)
frame_vm_group_bin_9335 = frame (4k)
frame_vm_group_bin_9336 = frame (4k)
frame_vm_group_bin_9337 = frame (4k)
frame_vm_group_bin_9338 = frame (4k)
frame_vm_group_bin_9339 = frame (4k)
frame_vm_group_bin_9340 = frame (4k)
frame_vm_group_bin_9341 = frame (4k)
frame_vm_group_bin_9342 = frame (4k)
frame_vm_group_bin_9343 = frame (4k)
frame_vm_group_bin_9344 = frame (4k)
frame_vm_group_bin_9345 = frame (4k)
frame_vm_group_bin_9346 = frame (4k)
frame_vm_group_bin_9347 = frame (4k)
frame_vm_group_bin_9348 = frame (4k)
frame_vm_group_bin_9349 = frame (4k)
frame_vm_group_bin_9350 = frame (4k)
frame_vm_group_bin_9351 = frame (4k)
frame_vm_group_bin_9352 = frame (4k)
frame_vm_group_bin_9353 = frame (4k)
frame_vm_group_bin_9354 = frame (4k)
frame_vm_group_bin_9355 = frame (4k)
frame_vm_group_bin_9356 = frame (4k)
frame_vm_group_bin_9357 = frame (4k)
frame_vm_group_bin_9358 = frame (4k)
frame_vm_group_bin_9359 = frame (4k)
frame_vm_group_bin_9360 = frame (4k)
frame_vm_group_bin_9361 = frame (4k)
frame_vm_group_bin_9362 = frame (4k)
frame_vm_group_bin_9363 = frame (4k)
frame_vm_group_bin_9364 = frame (4k)
frame_vm_group_bin_9365 = frame (4k)
frame_vm_group_bin_9366 = frame (4k)
frame_vm_group_bin_9367 = frame (4k)
frame_vm_group_bin_9368 = frame (4k)
frame_vm_group_bin_9369 = frame (4k)
frame_vm_group_bin_9370 = frame (4k)
frame_vm_group_bin_9371 = frame (4k)
frame_vm_group_bin_9372 = frame (4k)
frame_vm_group_bin_9373 = frame (4k)
frame_vm_group_bin_9374 = frame (4k)
frame_vm_group_bin_9375 = frame (4k)
frame_vm_group_bin_9376 = frame (4k)
frame_vm_group_bin_9377 = frame (4k)
frame_vm_group_bin_9378 = frame (4k)
frame_vm_group_bin_9379 = frame (4k)
frame_vm_group_bin_9380 = frame (4k)
frame_vm_group_bin_9381 = frame (4k)
frame_vm_group_bin_9382 = frame (4k)
frame_vm_group_bin_9383 = frame (4k)
frame_vm_group_bin_9384 = frame (4k)
frame_vm_group_bin_9385 = frame (4k)
frame_vm_group_bin_9386 = frame (4k)
frame_vm_group_bin_9387 = frame (4k)
frame_vm_group_bin_9388 = frame (4k)
frame_vm_group_bin_9389 = frame (4k)
frame_vm_group_bin_9390 = frame (4k)
frame_vm_group_bin_9391 = frame (4k)
frame_vm_group_bin_9392 = frame (4k)
frame_vm_group_bin_9393 = frame (4k)
frame_vm_group_bin_9394 = frame (4k)
frame_vm_group_bin_9395 = frame (4k)
frame_vm_group_bin_9396 = frame (4k)
frame_vm_group_bin_9397 = frame (4k)
frame_vm_group_bin_9398 = frame (4k)
frame_vm_group_bin_9399 = frame (4k)
frame_vm_group_bin_9400 = frame (4k)
frame_vm_group_bin_9401 = frame (4k)
frame_vm_group_bin_9402 = frame (4k)
frame_vm_group_bin_9403 = frame (4k)
frame_vm_group_bin_9404 = frame (4k)
frame_vm_group_bin_9405 = frame (4k)
frame_vm_group_bin_9406 = frame (4k)
frame_vm_group_bin_9407 = frame (4k)
frame_vm_group_bin_9408 = frame (4k)
frame_vm_group_bin_9409 = frame (4k)
frame_vm_group_bin_9410 = frame (4k)
frame_vm_group_bin_9411 = frame (4k)
frame_vm_group_bin_9412 = frame (4k)
frame_vm_group_bin_9413 = frame (4k)
frame_vm_group_bin_9414 = frame (4k)
frame_vm_group_bin_9415 = frame (4k)
frame_vm_group_bin_9416 = frame (4k)
frame_vm_group_bin_9417 = frame (4k)
frame_vm_group_bin_9418 = frame (4k)
frame_vm_group_bin_9419 = frame (4k)
frame_vm_group_bin_9420 = frame (4k)
frame_vm_group_bin_9421 = frame (4k)
frame_vm_group_bin_9422 = frame (4k)
frame_vm_group_bin_9423 = frame (4k)
frame_vm_group_bin_9424 = frame (4k)
frame_vm_group_bin_9425 = frame (4k)
frame_vm_group_bin_9426 = frame (4k)
frame_vm_group_bin_9427 = frame (4k)
frame_vm_group_bin_9428 = frame (4k)
frame_vm_group_bin_9429 = frame (4k)
frame_vm_group_bin_9430 = frame (4k)
frame_vm_group_bin_9431 = frame (4k)
frame_vm_group_bin_9432 = frame (4k)
frame_vm_group_bin_9433 = frame (4k)
frame_vm_group_bin_9434 = frame (4k)
frame_vm_group_bin_9435 = frame (4k)
frame_vm_group_bin_9436 = frame (4k)
frame_vm_group_bin_9437 = frame (4k)
frame_vm_group_bin_9438 = frame (4k)
frame_vm_group_bin_9439 = frame (4k)
frame_vm_group_bin_9440 = frame (4k)
frame_vm_group_bin_9441 = frame (4k)
frame_vm_group_bin_9442 = frame (4k)
frame_vm_group_bin_9443 = frame (4k)
frame_vm_group_bin_9444 = frame (4k)
frame_vm_group_bin_9445 = frame (4k)
frame_vm_group_bin_9446 = frame (4k)
frame_vm_group_bin_9447 = frame (4k)
frame_vm_group_bin_9448 = frame (4k)
frame_vm_group_bin_9449 = frame (4k)
frame_vm_group_bin_9450 = frame (4k)
frame_vm_group_bin_9451 = frame (4k)
frame_vm_group_bin_9452 = frame (4k)
frame_vm_group_bin_9453 = frame (4k)
frame_vm_group_bin_9454 = frame (4k)
frame_vm_group_bin_9455 = frame (4k)
frame_vm_group_bin_9456 = frame (4k)
frame_vm_group_bin_9457 = frame (4k)
frame_vm_group_bin_9458 = frame (4k)
frame_vm_group_bin_9459 = frame (4k)
frame_vm_group_bin_9460 = frame (4k)
frame_vm_group_bin_9461 = frame (4k)
frame_vm_group_bin_9462 = frame (4k)
frame_vm_group_bin_9463 = frame (4k)
frame_vm_group_bin_9464 = frame (4k)
frame_vm_group_bin_9465 = frame (4k)
frame_vm_group_bin_9466 = frame (4k)
frame_vm_group_bin_9467 = frame (4k)
frame_vm_group_bin_9468 = frame (4k)
frame_vm_group_bin_9469 = frame (4k)
frame_vm_group_bin_9470 = frame (4k)
frame_vm_group_bin_9471 = frame (4k)
frame_vm_group_bin_9472 = frame (4k)
frame_vm_group_bin_9473 = frame (4k)
frame_vm_group_bin_9474 = frame (4k)
frame_vm_group_bin_9475 = frame (4k)
frame_vm_group_bin_9476 = frame (4k)
frame_vm_group_bin_9477 = frame (4k)
frame_vm_group_bin_9478 = frame (4k)
frame_vm_group_bin_9479 = frame (4k)
frame_vm_group_bin_9480 = frame (4k)
frame_vm_group_bin_9481 = frame (4k)
frame_vm_group_bin_9482 = frame (4k)
frame_vm_group_bin_9483 = frame (4k)
frame_vm_group_bin_9484 = frame (4k)
frame_vm_group_bin_9485 = frame (4k)
frame_vm_group_bin_9486 = frame (4k)
frame_vm_group_bin_9487 = frame (4k)
frame_vm_group_bin_9488 = frame (4k)
frame_vm_group_bin_9489 = frame (4k)
frame_vm_group_bin_9490 = frame (4k)
frame_vm_group_bin_9491 = frame (4k)
frame_vm_group_bin_9492 = frame (4k)
frame_vm_group_bin_9493 = frame (4k)
frame_vm_group_bin_9494 = frame (4k)
frame_vm_group_bin_9495 = frame (4k)
frame_vm_group_bin_9496 = frame (4k)
frame_vm_group_bin_9497 = frame (4k)
frame_vm_group_bin_9498 = frame (4k)
frame_vm_group_bin_9499 = frame (4k)
frame_vm_group_bin_9500 = frame (4k)
frame_vm_group_bin_9501 = frame (4k)
frame_vm_group_bin_9502 = frame (4k)
frame_vm_group_bin_9503 = frame (4k)
frame_vm_group_bin_9504 = frame (4k)
frame_vm_group_bin_9505 = frame (4k)
frame_vm_group_bin_9506 = frame (4k)
frame_vm_group_bin_9507 = frame (4k)
frame_vm_group_bin_9508 = frame (4k)
frame_vm_group_bin_9509 = frame (4k)
frame_vm_group_bin_9510 = frame (4k)
frame_vm_group_bin_9511 = frame (4k)
frame_vm_group_bin_9512 = frame (4k)
frame_vm_group_bin_9513 = frame (4k)
frame_vm_group_bin_9514 = frame (4k)
frame_vm_group_bin_9515 = frame (4k)
frame_vm_group_bin_9516 = frame (4k)
frame_vm_group_bin_9517 = frame (4k)
frame_vm_group_bin_9518 = frame (4k)
frame_vm_group_bin_9519 = frame (4k)
frame_vm_group_bin_9520 = frame (4k)
frame_vm_group_bin_9521 = frame (4k)
frame_vm_group_bin_9522 = frame (4k)
frame_vm_group_bin_9523 = frame (4k)
frame_vm_group_bin_9524 = frame (4k)
frame_vm_group_bin_9525 = frame (4k)
frame_vm_group_bin_9526 = frame (4k)
frame_vm_group_bin_9527 = frame (4k)
frame_vm_group_bin_9528 = frame (4k)
frame_vm_group_bin_9529 = frame (4k)
frame_vm_group_bin_9530 = frame (4k)
frame_vm_group_bin_9531 = frame (4k)
frame_vm_group_bin_9532 = frame (4k)
frame_vm_group_bin_9533 = frame (4k)
frame_vm_group_bin_9534 = frame (4k)
frame_vm_group_bin_9535 = frame (4k)
frame_vm_group_bin_9536 = frame (4k)
frame_vm_group_bin_9537 = frame (4k)
frame_vm_group_bin_9538 = frame (4k)
frame_vm_group_bin_9539 = frame (4k)
frame_vm_group_bin_9540 = frame (4k)
frame_vm_group_bin_9541 = frame (4k)
frame_vm_group_bin_9542 = frame (4k)
frame_vm_group_bin_9543 = frame (4k)
frame_vm_group_bin_9544 = frame (4k)
frame_vm_group_bin_9545 = frame (4k)
frame_vm_group_bin_9546 = frame (4k)
frame_vm_group_bin_9547 = frame (4k)
frame_vm_group_bin_9548 = frame (4k)
frame_vm_group_bin_9549 = frame (4k)
frame_vm_group_bin_9550 = frame (4k)
frame_vm_group_bin_9551 = frame (4k)
frame_vm_group_bin_9552 = frame (4k)
frame_vm_group_bin_9553 = frame (4k)
frame_vm_group_bin_9554 = frame (4k)
frame_vm_group_bin_9555 = frame (4k)
frame_vm_group_bin_9556 = frame (4k)
frame_vm_group_bin_9557 = frame (4k)
frame_vm_group_bin_9558 = frame (4k)
frame_vm_group_bin_9559 = frame (4k)
frame_vm_group_bin_9560 = frame (4k)
frame_vm_group_bin_9561 = frame (4k)
frame_vm_group_bin_9562 = frame (4k)
frame_vm_group_bin_9563 = frame (4k)
frame_vm_group_bin_9564 = frame (4k)
frame_vm_group_bin_9565 = frame (4k)
frame_vm_group_bin_9566 = frame (4k)
frame_vm_group_bin_9567 = frame (4k)
frame_vm_group_bin_9568 = frame (4k)
frame_vm_group_bin_9569 = frame (4k)
frame_vm_group_bin_9570 = frame (4k)
frame_vm_group_bin_9571 = frame (4k)
frame_vm_group_bin_9572 = frame (4k)
frame_vm_group_bin_9573 = frame (4k)
frame_vm_group_bin_9574 = frame (4k)
frame_vm_group_bin_9575 = frame (4k)
frame_vm_group_bin_9576 = frame (4k)
frame_vm_group_bin_9577 = frame (4k)
frame_vm_group_bin_9578 = frame (4k)
frame_vm_group_bin_9579 = frame (4k)
frame_vm_group_bin_9580 = frame (4k)
frame_vm_group_bin_9581 = frame (4k)
frame_vm_group_bin_9582 = frame (4k)
frame_vm_group_bin_9583 = frame (4k)
frame_vm_group_bin_9584 = frame (4k)
frame_vm_group_bin_9585 = frame (4k)
frame_vm_group_bin_9586 = frame (4k)
frame_vm_group_bin_9587 = frame (4k)
frame_vm_group_bin_9588 = frame (4k)
frame_vm_group_bin_9589 = frame (4k)
frame_vm_group_bin_9590 = frame (4k)
frame_vm_group_bin_9591 = frame (4k)
frame_vm_group_bin_9592 = frame (4k)
frame_vm_group_bin_9593 = frame (4k)
frame_vm_group_bin_9594 = frame (4k)
frame_vm_group_bin_9595 = frame (4k)
frame_vm_group_bin_9596 = frame (4k)
frame_vm_group_bin_9597 = frame (4k)
frame_vm_group_bin_9598 = frame (4k)
frame_vm_group_bin_9599 = frame (4k)
frame_vm_group_bin_9600 = frame (4k)
frame_vm_group_bin_9601 = frame (4k)
frame_vm_group_bin_9602 = frame (4k)
frame_vm_group_bin_9603 = frame (4k)
frame_vm_group_bin_9604 = frame (4k)
frame_vm_group_bin_9605 = frame (4k)
frame_vm_group_bin_9606 = frame (4k)
frame_vm_group_bin_9607 = frame (4k)
frame_vm_group_bin_9608 = frame (4k)
frame_vm_group_bin_9609 = frame (4k)
frame_vm_group_bin_9610 = frame (4k)
frame_vm_group_bin_9611 = frame (4k)
frame_vm_group_bin_9612 = frame (4k)
frame_vm_group_bin_9613 = frame (4k)
frame_vm_group_bin_9614 = frame (4k)
frame_vm_group_bin_9615 = frame (4k)
frame_vm_group_bin_9616 = frame (4k)
frame_vm_group_bin_9617 = frame (4k)
frame_vm_group_bin_9618 = frame (4k)
frame_vm_group_bin_9619 = frame (4k)
frame_vm_group_bin_9620 = frame (4k)
frame_vm_group_bin_9621 = frame (4k)
frame_vm_group_bin_9622 = frame (4k)
frame_vm_group_bin_9623 = frame (4k)
frame_vm_group_bin_9624 = frame (4k)
frame_vm_group_bin_9625 = frame (4k)
frame_vm_group_bin_9626 = frame (4k)
frame_vm_group_bin_9627 = frame (4k)
frame_vm_group_bin_9628 = frame (4k)
frame_vm_group_bin_9629 = frame (4k)
frame_vm_group_bin_9630 = frame (4k)
frame_vm_group_bin_9631 = frame (4k)
frame_vm_group_bin_9632 = frame (4k)
frame_vm_group_bin_9633 = frame (4k)
frame_vm_group_bin_9634 = frame (4k)
frame_vm_group_bin_9635 = frame (4k)
frame_vm_group_bin_9636 = frame (4k)
frame_vm_group_bin_9637 = frame (4k)
frame_vm_group_bin_9638 = frame (4k)
frame_vm_group_bin_9639 = frame (4k)
frame_vm_group_bin_9640 = frame (4k)
frame_vm_group_bin_9641 = frame (4k)
frame_vm_group_bin_9642 = frame (4k)
frame_vm_group_bin_9643 = frame (4k)
frame_vm_group_bin_9644 = frame (4k)
frame_vm_group_bin_9645 = frame (4k)
frame_vm_group_bin_9646 = frame (4k)
frame_vm_group_bin_9647 = frame (4k)
frame_vm_group_bin_9648 = frame (4k)
frame_vm_group_bin_9649 = frame (4k)
frame_vm_group_bin_9650 = frame (4k)
frame_vm_group_bin_9651 = frame (4k)
frame_vm_group_bin_9652 = frame (4k)
frame_vm_group_bin_9653 = frame (4k)
frame_vm_group_bin_9654 = frame (4k)
frame_vm_group_bin_9655 = frame (4k)
frame_vm_group_bin_9656 = frame (4k)
frame_vm_group_bin_9657 = frame (4k)
frame_vm_group_bin_9658 = frame (4k)
frame_vm_group_bin_9659 = frame (4k)
frame_vm_group_bin_9660 = frame (4k)
frame_vm_group_bin_9661 = frame (4k)
frame_vm_group_bin_9662 = frame (4k)
frame_vm_group_bin_9663 = frame (4k)
frame_vm_group_bin_9664 = frame (4k)
frame_vm_group_bin_9665 = frame (4k)
frame_vm_group_bin_9666 = frame (4k)
frame_vm_group_bin_9667 = frame (4k)
frame_vm_group_bin_9668 = frame (4k)
frame_vm_group_bin_9669 = frame (4k)
frame_vm_group_bin_9670 = frame (4k)
frame_vm_group_bin_9671 = frame (4k)
frame_vm_group_bin_9672 = frame (4k)
frame_vm_group_bin_9673 = frame (4k)
frame_vm_group_bin_9674 = frame (4k)
frame_vm_group_bin_9675 = frame (4k)
frame_vm_group_bin_9676 = frame (4k)
frame_vm_group_bin_9677 = frame (4k)
frame_vm_group_bin_9678 = frame (4k)
frame_vm_group_bin_9679 = frame (4k)
frame_vm_group_bin_9680 = frame (4k)
frame_vm_group_bin_9681 = frame (4k)
frame_vm_group_bin_9682 = frame (4k)
frame_vm_group_bin_9683 = frame (4k)
frame_vm_group_bin_9684 = frame (4k)
frame_vm_group_bin_9685 = frame (4k)
frame_vm_group_bin_9686 = frame (4k)
frame_vm_group_bin_9687 = frame (4k)
frame_vm_group_bin_9688 = frame (4k)
frame_vm_group_bin_9689 = frame (4k)
frame_vm_group_bin_9690 = frame (4k)
frame_vm_group_bin_9691 = frame (4k)
frame_vm_group_bin_9692 = frame (4k)
frame_vm_group_bin_9693 = frame (4k)
frame_vm_group_bin_9694 = frame (4k)
frame_vm_group_bin_9695 = frame (4k)
frame_vm_group_bin_9696 = frame (4k)
frame_vm_group_bin_9697 = frame (4k)
frame_vm_group_bin_9698 = frame (4k)
frame_vm_group_bin_9699 = frame (4k)
frame_vm_group_bin_9700 = frame (4k)
frame_vm_group_bin_9701 = frame (4k)
frame_vm_group_bin_9702 = frame (4k)
frame_vm_group_bin_9703 = frame (4k)
frame_vm_group_bin_9704 = frame (4k)
frame_vm_group_bin_9705 = frame (4k)
frame_vm_group_bin_9706 = frame (4k)
frame_vm_group_bin_9707 = frame (4k)
frame_vm_group_bin_9708 = frame (4k)
frame_vm_group_bin_9709 = frame (4k)
frame_vm_group_bin_9710 = frame (4k)
frame_vm_group_bin_9711 = frame (4k)
frame_vm_group_bin_9712 = frame (4k)
frame_vm_group_bin_9713 = frame (4k)
frame_vm_group_bin_9714 = frame (4k)
frame_vm_group_bin_9715 = frame (4k)
frame_vm_group_bin_9716 = frame (4k)
frame_vm_group_bin_9717 = frame (4k)
frame_vm_group_bin_9718 = frame (4k)
frame_vm_group_bin_9719 = frame (4k)
frame_vm_group_bin_9720 = frame (4k)
frame_vm_group_bin_9721 = frame (4k)
frame_vm_group_bin_9722 = frame (4k)
frame_vm_group_bin_9723 = frame (4k)
frame_vm_group_bin_9724 = frame (4k)
frame_vm_group_bin_9725 = frame (4k)
frame_vm_group_bin_9726 = frame (4k)
frame_vm_group_bin_9727 = frame (4k)
frame_vm_group_bin_9728 = frame (4k)
frame_vm_group_bin_9729 = frame (4k)
frame_vm_group_bin_9730 = frame (4k)
frame_vm_group_bin_9731 = frame (4k)
frame_vm_group_bin_9732 = frame (4k)
frame_vm_group_bin_9733 = frame (4k)
frame_vm_group_bin_9734 = frame (4k)
frame_vm_group_bin_9735 = frame (4k)
frame_vm_group_bin_9736 = frame (4k)
frame_vm_group_bin_9737 = frame (4k)
frame_vm_group_bin_9738 = frame (4k)
frame_vm_group_bin_9739 = frame (4k)
frame_vm_group_bin_9740 = frame (4k)
frame_vm_group_bin_9741 = frame (4k)
frame_vm_group_bin_9742 = frame (4k)
frame_vm_group_bin_9743 = frame (4k)
frame_vm_group_bin_9744 = frame (4k)
frame_vm_group_bin_9745 = frame (4k)
frame_vm_group_bin_9746 = frame (4k)
frame_vm_group_bin_9747 = frame (4k)
frame_vm_group_bin_9748 = frame (4k)
frame_vm_group_bin_9749 = frame (4k)
frame_vm_group_bin_9750 = frame (4k)
frame_vm_group_bin_9751 = frame (4k)
frame_vm_group_bin_9752 = frame (4k)
frame_vm_group_bin_9753 = frame (4k)
frame_vm_group_bin_9754 = frame (4k)
frame_vm_group_bin_9755 = frame (4k)
frame_vm_group_bin_9756 = frame (4k)
frame_vm_group_bin_9757 = frame (4k)
frame_vm_group_bin_9758 = frame (4k)
frame_vm_group_bin_9759 = frame (4k)
frame_vm_group_bin_9760 = frame (4k)
frame_vm_group_bin_9761 = frame (4k)
frame_vm_group_bin_9762 = frame (4k)
frame_vm_group_bin_9763 = frame (4k)
frame_vm_group_bin_9764 = frame (4k)
frame_vm_group_bin_9765 = frame (4k)
frame_vm_group_bin_9766 = frame (4k)
frame_vm_group_bin_9767 = frame (4k)
frame_vm_group_bin_9768 = frame (4k)
frame_vm_group_bin_9769 = frame (4k)
frame_vm_group_bin_9770 = frame (4k)
frame_vm_group_bin_9771 = frame (4k)
frame_vm_group_bin_9772 = frame (4k)
frame_vm_group_bin_9773 = frame (4k)
frame_vm_group_bin_9774 = frame (4k)
frame_vm_group_bin_9775 = frame (4k)
frame_vm_group_bin_9776 = frame (4k)
frame_vm_group_bin_9777 = frame (4k)
frame_vm_group_bin_9778 = frame (4k)
frame_vm_group_bin_9779 = frame (4k)
frame_vm_group_bin_9780 = frame (4k)
frame_vm_group_bin_9781 = frame (4k)
frame_vm_group_bin_9782 = frame (4k)
frame_vm_group_bin_9783 = frame (4k)
frame_vm_group_bin_9784 = frame (4k)
frame_vm_group_bin_9785 = frame (4k)
frame_vm_group_bin_9786 = frame (4k)
frame_vm_group_bin_9787 = frame (4k)
frame_vm_group_bin_9788 = frame (4k)
frame_vm_group_bin_9789 = frame (4k)
frame_vm_group_bin_9790 = frame (4k)
frame_vm_group_bin_9791 = frame (4k)
frame_vm_group_bin_9792 = frame (4k)
frame_vm_group_bin_9793 = frame (4k)
frame_vm_group_bin_9794 = frame (4k)
frame_vm_group_bin_9795 = frame (4k)
frame_vm_group_bin_9796 = frame (4k)
frame_vm_group_bin_9797 = frame (4k)
frame_vm_group_bin_9798 = frame (4k)
frame_vm_group_bin_9799 = frame (4k)
frame_vm_group_bin_9800 = frame (4k)
frame_vm_group_bin_9801 = frame (4k)
frame_vm_group_bin_9802 = frame (4k)
frame_vm_group_bin_9803 = frame (4k)
frame_vm_group_bin_9804 = frame (4k)
frame_vm_group_bin_9805 = frame (4k)
frame_vm_group_bin_9806 = frame (4k)
frame_vm_group_bin_9807 = frame (4k)
frame_vm_group_bin_9808 = frame (4k)
frame_vm_group_bin_9809 = frame (4k)
frame_vm_group_bin_9810 = frame (4k)
frame_vm_group_bin_9811 = frame (4k)
frame_vm_group_bin_9812 = frame (4k)
frame_vm_group_bin_9813 = frame (4k)
frame_vm_group_bin_9814 = frame (4k)
frame_vm_group_bin_9815 = frame (4k)
frame_vm_group_bin_9816 = frame (4k)
frame_vm_group_bin_9817 = frame (4k)
frame_vm_group_bin_9818 = frame (4k)
frame_vm_group_bin_9819 = frame (4k)
frame_vm_group_bin_9820 = frame (4k)
frame_vm_group_bin_9821 = frame (4k)
frame_vm_group_bin_9822 = frame (4k)
frame_vm_group_bin_9823 = frame (4k)
frame_vm_group_bin_9824 = frame (4k)
frame_vm_group_bin_9825 = frame (4k)
frame_vm_group_bin_9826 = frame (4k)
frame_vm_group_bin_9827 = frame (4k)
frame_vm_group_bin_9828 = frame (4k)
frame_vm_group_bin_9829 = frame (4k)
frame_vm_group_bin_9830 = frame (4k)
frame_vm_group_bin_9831 = frame (4k)
frame_vm_group_bin_9832 = frame (4k)
frame_vm_group_bin_9833 = frame (4k)
frame_vm_group_bin_9834 = frame (4k)
frame_vm_group_bin_9835 = frame (4k)
frame_vm_group_bin_9836 = frame (4k)
frame_vm_group_bin_9837 = frame (4k)
frame_vm_group_bin_9838 = frame (4k)
frame_vm_group_bin_9839 = frame (4k)
frame_vm_group_bin_9840 = frame (4k)
frame_vm_group_bin_9841 = frame (4k)
frame_vm_group_bin_9842 = frame (4k)
frame_vm_group_bin_9843 = frame (4k)
frame_vm_group_bin_9844 = frame (4k)
frame_vm_group_bin_9845 = frame (4k)
frame_vm_group_bin_9846 = frame (4k)
frame_vm_group_bin_9847 = frame (4k)
frame_vm_group_bin_9848 = frame (4k)
frame_vm_group_bin_9849 = frame (4k)
frame_vm_group_bin_9850 = frame (4k)
frame_vm_group_bin_9851 = frame (4k)
frame_vm_group_bin_9852 = frame (4k)
frame_vm_group_bin_9853 = frame (4k)
frame_vm_group_bin_9854 = frame (4k)
frame_vm_group_bin_9855 = frame (4k)
frame_vm_group_bin_9856 = frame (4k)
frame_vm_group_bin_9857 = frame (4k)
frame_vm_group_bin_9858 = frame (4k)
frame_vm_group_bin_9859 = frame (4k)
frame_vm_group_bin_9860 = frame (4k)
frame_vm_group_bin_9861 = frame (4k)
frame_vm_group_bin_9862 = frame (4k)
frame_vm_group_bin_9863 = frame (4k)
frame_vm_group_bin_9864 = frame (4k)
frame_vm_group_bin_9865 = frame (4k)
frame_vm_group_bin_9866 = frame (4k)
frame_vm_group_bin_9867 = frame (4k)
frame_vm_group_bin_9868 = frame (4k)
frame_vm_group_bin_9869 = frame (4k)
frame_vm_group_bin_9870 = frame (4k)
frame_vm_group_bin_9871 = frame (4k)
frame_vm_group_bin_9872 = frame (4k)
frame_vm_group_bin_9873 = frame (4k)
frame_vm_group_bin_9874 = frame (4k)
frame_vm_group_bin_9875 = frame (4k)
frame_vm_group_bin_9876 = frame (4k)
frame_vm_group_bin_9877 = frame (4k)
frame_vm_group_bin_9878 = frame (4k)
frame_vm_group_bin_9879 = frame (4k)
frame_vm_group_bin_9880 = frame (4k)
frame_vm_group_bin_9881 = frame (4k)
frame_vm_group_bin_9882 = frame (4k)
frame_vm_group_bin_9883 = frame (4k)
frame_vm_group_bin_9884 = frame (4k)
frame_vm_group_bin_9885 = frame (4k)
frame_vm_group_bin_9886 = frame (4k)
frame_vm_group_bin_9887 = frame (4k)
frame_vm_group_bin_9888 = frame (4k)
frame_vm_group_bin_9889 = frame (4k)
frame_vm_group_bin_9890 = frame (4k)
frame_vm_group_bin_9891 = frame (4k)
frame_vm_group_bin_9892 = frame (4k)
frame_vm_group_bin_9893 = frame (4k)
frame_vm_group_bin_9894 = frame (4k)
frame_vm_group_bin_9895 = frame (4k)
frame_vm_group_bin_9896 = frame (4k)
frame_vm_group_bin_9897 = frame (4k)
frame_vm_group_bin_9898 = frame (4k)
frame_vm_group_bin_9899 = frame (4k)
frame_vm_group_bin_9900 = frame (4k)
frame_vm_group_bin_9901 = frame (4k)
frame_vm_group_bin_9902 = frame (4k)
frame_vm_group_bin_9903 = frame (4k)
frame_vm_group_bin_9904 = frame (4k)
frame_vm_group_bin_9905 = frame (4k)
frame_vm_group_bin_9906 = frame (4k)
frame_vm_group_bin_9907 = frame (4k)
frame_vm_group_bin_9908 = frame (4k)
frame_vm_group_bin_9909 = frame (4k)
frame_vm_group_bin_9910 = frame (4k)
frame_vm_group_bin_9911 = frame (4k)
frame_vm_group_bin_9912 = frame (4k)
frame_vm_group_bin_9913 = frame (4k)
frame_vm_group_bin_9914 = frame (4k)
frame_vm_group_bin_9915 = frame (4k)
frame_vm_group_bin_9916 = frame (4k)
frame_vm_group_bin_9917 = frame (4k)
frame_vm_group_bin_9918 = frame (4k)
frame_vm_group_bin_9919 = frame (4k)
frame_vm_group_bin_9920 = frame (4k)
frame_vm_group_bin_9921 = frame (4k)
frame_vm_group_bin_9922 = frame (4k)
frame_vm_group_bin_9923 = frame (4k)
frame_vm_group_bin_9924 = frame (4k)
frame_vm_group_bin_9925 = frame (4k)
frame_vm_group_bin_9926 = frame (4k)
frame_vm_group_bin_9927 = frame (4k)
frame_vm_group_bin_9928 = frame (4k)
frame_vm_group_bin_9929 = frame (4k)
frame_vm_group_bin_9930 = frame (4k)
frame_vm_group_bin_9931 = frame (4k)
frame_vm_group_bin_9932 = frame (4k)
frame_vm_group_bin_9933 = frame (4k)
frame_vm_group_bin_9934 = frame (4k)
frame_vm_group_bin_9935 = frame (4k)
frame_vm_group_bin_9936 = frame (4k)
frame_vm_group_bin_9937 = frame (4k)
frame_vm_group_bin_9938 = frame (4k)
frame_vm_group_bin_9939 = frame (4k)
frame_vm_group_bin_9940 = frame (4k)
frame_vm_group_bin_9941 = frame (4k)
frame_vm_group_bin_9942 = frame (4k)
frame_vm_group_bin_9943 = frame (4k)
frame_vm_group_bin_9944 = frame (4k)
frame_vm_group_bin_9945 = frame (4k)
frame_vm_group_bin_9946 = frame (4k)
frame_vm_group_bin_9947 = frame (4k)
frame_vm_group_bin_9948 = frame (4k)
frame_vm_group_bin_9949 = frame (4k)
frame_vm_group_bin_9950 = frame (4k)
frame_vm_group_bin_9951 = frame (4k)
frame_vm_group_bin_9952 = frame (4k)
frame_vm_group_bin_9953 = frame (4k)
frame_vm_group_bin_9954 = frame (4k)
frame_vm_group_bin_9955 = frame (4k)
frame_vm_group_bin_9956 = frame (4k)
frame_vm_group_bin_9957 = frame (4k)
frame_vm_group_bin_9958 = frame (4k)
frame_vm_group_bin_9959 = frame (4k)
frame_vm_group_bin_9960 = frame (4k)
frame_vm_group_bin_9961 = frame (4k)
frame_vm_group_bin_9962 = frame (4k)
frame_vm_group_bin_9963 = frame (4k)
frame_vm_group_bin_9964 = frame (4k)
frame_vm_group_bin_9965 = frame (4k)
frame_vm_group_bin_9966 = frame (4k)
frame_vm_group_bin_9967 = frame (4k)
frame_vm_group_bin_9968 = frame (4k)
frame_vm_group_bin_9969 = frame (4k)
frame_vm_group_bin_9970 = frame (4k)
frame_vm_group_bin_9971 = frame (4k)
frame_vm_group_bin_9972 = frame (4k)
frame_vm_group_bin_9973 = frame (4k)
frame_vm_group_bin_9974 = frame (4k)
frame_vm_group_bin_9975 = frame (4k)
frame_vm_group_bin_9976 = frame (4k)
frame_vm_group_bin_9977 = frame (4k)
frame_vm_group_bin_9978 = frame (4k)
frame_vm_group_bin_9979 = frame (4k)
frame_vm_group_bin_9980 = frame (4k)
frame_vm_group_bin_9981 = frame (4k)
frame_vm_group_bin_9982 = frame (4k)
frame_vm_group_bin_9983 = frame (4k)
frame_vm_group_bin_9984 = frame (4k)
frame_vm_group_bin_9985 = frame (4k)
frame_vm_group_bin_9986 = frame (4k)
frame_vm_group_bin_9987 = frame (4k)
frame_vm_group_bin_9988 = frame (4k)
frame_vm_group_bin_9989 = frame (4k)
frame_vm_group_bin_9990 = frame (4k)
frame_vm_group_bin_9991 = frame (4k)
frame_vm_group_bin_9992 = frame (4k)
frame_vm_group_bin_9993 = frame (4k)
frame_vm_group_bin_9994 = frame (4k)
frame_vm_group_bin_9995 = frame (4k)
frame_vm_group_bin_9996 = frame (4k)
frame_vm_group_bin_9997 = frame (4k)
frame_vm_group_bin_9998 = frame (4k)
frame_vm_group_bin_9999 = frame (4k)
gcs_recv_inf.px4_recv_inf_ep = ep
gpio_can_intAck_handoff_0 = ep
gpio_can_intAck_lock_0 = notification
gpio_can_intAck_notification_0 = notification
gpio_can_int_handoff_0 = ep
gpio_can_int_lock_0 = notification
gpio_can_int_notification_0 = notification
gpio_grp26_irq_irq = irq
gpio_grp26_irq_ntfn = notification
gpio_grp28_irq_irq = irq
gpio_grp28_irq_ntfn = notification
gpio_grp31_irq_irq = irq
gpio_grp31_irq_ntfn = notification
gpio_obj_8_0_control_9_tcb = tcb (addr: 0x14de00, ip: 0x18af0, sp: 0x17e000, elf: gpio_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [1], fault_ep: 0x00000002)
gpio_obj_8_0_fault_handler_15_0000_tcb = tcb (addr: 0x138e00, ip: 0x18af0, sp: 0x154000, elf: gpio_obj_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [15])
gpio_obj_8_CANIntAck_9_0000_tcb = tcb (addr: 0x13be00, ip: 0x18af0, sp: 0x15a000, elf: gpio_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [13], fault_ep: 0x0000000e)
gpio_obj_8_gpio_4_0000_tcb = tcb (addr: 0x13ee00, ip: 0x18af0, sp: 0x160000, elf: gpio_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [11], fault_ep: 0x0000000c)
gpio_obj_8_irq_grp26_int_13_0000_tcb = tcb (addr: 0x147e00, ip: 0x18af0, sp: 0x172000, elf: gpio_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [5], fault_ep: 0x00000006)
gpio_obj_8_irq_grp28_int_13_0000_tcb = tcb (addr: 0x14ae00, ip: 0x18af0, sp: 0x178000, elf: gpio_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [3], fault_ep: 0x00000004)
gpio_obj_8_irq_grp31_int_13_0000_tcb = tcb (addr: 0x144e00, ip: 0x18af0, sp: 0x16c000, elf: gpio_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [7], fault_ep: 0x00000008)
gpio_obj_8_xint16_31_int_13_0000_tcb = tcb (addr: 0x141e00, ip: 0x18af0, sp: 0x166000, elf: gpio_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [9], fault_ep: 0x0000000a)
gpio_obj_cnode = cnode (6 bits)
gpio_obj_fault_ep = ep
gpio_obj_group_bin_pd = pd
gpio_obj_interface_init_ep = ep
gpio_obj_post_init_ep = ep
gpio_obj_pre_init_ep = ep
gpio_xint16_31_irq_irq = irq
gpio_xint16_31_irq_ntfn = notification
i2c0_irq_irq = irq
i2c0_irq_ntfn = notification
pilot_obj_9_0_control_9_tcb = tcb (addr: 0x145e00, ip: 0x1a81c, sp: 0x158000, elf: pilot_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [1], fault_ep: 0x00000002)
pilot_obj_9_0_fault_handler_15_0000_tcb = tcb (addr: 0x13fe00, ip: 0x1a81c, sp: 0x14c000, elf: pilot_obj_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [5])
pilot_obj_9_mavlink_7_0000_tcb = tcb (addr: 0x142e00, ip: 0x1a81c, sp: 0x152000, elf: pilot_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [3], fault_ep: 0x00000004)
pilot_obj_cnode = cnode (5 bits)
pilot_obj_fault_ep = ep
pilot_obj_group_bin_pd = pd
pilot_obj_interface_init_ep = ep
pilot_obj_post_init_ep = ep
pilot_obj_pre_init_ep = ep
pt_can_obj_group_bin_0000 = pt
pt_clk_obj_group_bin_0000 = pt
pt_clk_obj_group_bin_0106 = pt
pt_clk_obj_group_bin_0285 = pt
pt_gpio_obj_group_bin_0000 = pt
pt_gpio_obj_group_bin_0007 = pt
pt_gpio_obj_group_bin_0052 = pt
pt_pilot_obj_group_bin_0000 = pt
pt_pwm_obj_group_bin_0000 = pt
pt_pwm_obj_group_bin_0259 = pt
pt_spi_obj_group_bin_0000 = pt
pt_spi_obj_group_bin_0247 = pt
pt_timer_obj_group_bin_0000 = pt
pt_timer_obj_group_bin_0235 = pt
pt_uart_gcs_group_bin_0000 = pt
pt_uart_gcs_group_bin_0246 = pt
pt_uart_px4_group_bin_0000 = pt
pt_uart_px4_group_bin_0246 = pt
pt_vm_group_bin_0000 = pt
pt_vm_group_bin_0002 = pt
pt_vm_group_bin_0004 = pt
pt_vm_group_bin_0006 = pt
pt_vm_group_bin_0008 = pt
pt_vm_group_bin_0010 = pt
pt_vm_group_bin_0012 = pt
pt_vm_group_bin_0014 = pt
pt_vm_group_bin_0016 = pt
pt_vm_group_bin_0018 = pt
pt_vm_group_bin_0020 = pt
pt_vm_group_bin_0022 = pt
pt_vm_group_bin_0024 = pt
pt_vm_group_bin_0026 = pt
pt_vm_group_bin_0028 = pt
pt_vm_group_bin_0031 = pt
pt_vm_group_bin_0033 = pt
pt_vm_group_bin_0035 = pt
pt_vm_group_bin_0037 = pt
pt_vm_group_bin_0039 = pt
pt_vm_group_bin_0044 = pt
pt_vm_group_bin_0051 = pt
pt_vm_group_bin_0054 = pt
pt_vm_group_bin_0060 = pt
pt_vm_group_bin_0063 = pt
pt_vm_group_bin_0065 = pt
pt_vm_group_bin_0071 = pt
pt_vm_group_bin_0079 = pt
pt_vm_group_bin_0099 = pt
pt_vm_group_bin_0107 = pt
pt_vm_group_bin_0115 = pt
pt_vm_group_bin_0117 = pt
pt_vm_group_bin_0123 = pt
pt_vm_group_bin_0134 = pt
pt_vm_group_bin_0167 = pt
pt_vm_group_bin_0176 = pt
pt_vm_group_bin_0196 = pt
pt_vm_group_bin_0203 = pt
pt_vm_group_bin_0210 = pt
pt_vm_group_bin_0220 = pt
pt_vm_group_bin_0239 = pt
pt_vm_group_bin_0272 = pt
pt_vm_group_bin_0328 = pt
pt_vm_group_bin_0380 = pt
pt_vm_group_bin_0403 = pt
pt_vm_group_bin_1120 = pt
pwm_obj_7_0_control_9_tcb = tcb (addr: 0x147e00, ip: 0x17b40, sp: 0x16c000, elf: pwm_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [4], fault_ep: 0x00000005)
pwm_obj_7_0_fault_handler_15_0000_tcb = tcb (addr: 0x138e00, ip: 0x17b40, sp: 0x14e000, elf: pwm_obj_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [14])
pwm_obj_7_i2c0_int_8_0000_tcb = tcb (addr: 0x144e00, ip: 0x17b40, sp: 0x166000, elf: pwm_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [6], fault_ep: 0x00000007)
pwm_obj_7_pwm_3_0000_tcb = tcb (addr: 0x13be00, ip: 0x17b40, sp: 0x154000, elf: pwm_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [12], fault_ep: 0x0000000d)
pwm_obj_7_signal_6_0000_tcb = tcb (addr: 0x141e00, ip: 0x17b40, sp: 0x160000, elf: pwm_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [8], fault_ep: 0x00000009)
pwm_obj_7_timer_update_12_0000_tcb = tcb (addr: 0x13ee00, ip: 0x17b40, sp: 0x15a000, elf: pwm_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [10], fault_ep: 0x0000000b)
pwm_obj_bus_sem = ep
pwm_obj_cnode = cnode (5 bits)
pwm_obj_fault_ep = ep
pwm_obj_group_bin_pd = pd
pwm_obj_interface_init_ep = ep
pwm_obj_post_init_ep = ep
pwm_obj_pre_init_ep = ep
pwm_obj_set_motors = notification
pwm_obj_sig = notification
pwm_sig_handoff_0 = ep
pwm_sig_lock_0 = notification
pwm_sig_notification_0 = notification
pwm_timer_handoff_0 = ep
pwm_timer_lock_0 = notification
pwm_timer_notification_0 = notification
restart_vm_handoff_0 = ep
restart_vm_lock_0 = notification
restart_vm_notification_0 = notification
spi1_irq_irq = irq
spi1_irq_ntfn = notification
spi_clk_ep = ep
spi_gpio_ep = ep
spi_obj_7_0_control_9_tcb = tcb (addr: 0x140e00, ip: 0x165bc, sp: 0x159000, elf: spi_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [2], fault_ep: 0x00000003)
spi_obj_7_0_fault_handler_15_0000_tcb = tcb (addr: 0x137e00, ip: 0x165bc, sp: 0x147000, elf: spi_obj_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [8])
spi_obj_7_spi1_int_8_0000_tcb = tcb (addr: 0x13de00, ip: 0x165bc, sp: 0x153000, elf: spi_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [4], fault_ep: 0x00000005)
spi_obj_7_spi_3_0000_tcb = tcb (addr: 0x13ae00, ip: 0x165bc, sp: 0x14d000, elf: spi_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [6], fault_ep: 0x00000007)
spi_obj_bus_sem = ep
spi_obj_cnode = cnode (5 bits)
spi_obj_fault_ep = ep
spi_obj_group_bin_pd = pd
spi_obj_interface_init_ep = ep
spi_obj_post_init_ep = ep
spi_obj_pre_init_ep = ep
timer_irq_irq = irq
timer_irq_ntfn = notification
timer_obj_9_0_control_9_tcb = tcb (addr: 0x137e00, ip: 0x14578, sp: 0x14a000, elf: timer_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [1], fault_ep: 0x00000002)
timer_obj_9_0_fault_handler_15_0000_tcb = tcb (addr: 0x131e00, ip: 0x14578, sp: 0x13e000, elf: timer_obj_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [5])
timer_obj_9_irq_3_0000_tcb = tcb (addr: 0x134e00, ip: 0x14578, sp: 0x144000, elf: timer_obj_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [3], fault_ep: 0x00000004)
timer_obj_cnode = cnode (4 bits)
timer_obj_fault_ep = ep
timer_obj_group_bin_pd = pd
timer_obj_interface_init_ep = ep
timer_obj_post_init_ep = ep
timer_obj_pre_init_ep = ep
uart_gcs_8_0_control_9_tcb = tcb (addr: 0x13de00, ip: 0x159b0, sp: 0x156000, elf: uart_gcs_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [3], fault_ep: 0x00000004)
uart_gcs_8_0_fault_handler_15_0000_tcb = tcb (addr: 0x134e00, ip: 0x159b0, sp: 0x144000, elf: uart_gcs_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [9])
uart_gcs_8_interrupt_9_0000_tcb = tcb (addr: 0x13ae00, ip: 0x159b0, sp: 0x150000, elf: uart_gcs_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [5], fault_ep: 0x00000006)
uart_gcs_8_uart_4_0000_tcb = tcb (addr: 0x137e00, ip: 0x159b0, sp: 0x14a000, elf: uart_gcs_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [7], fault_ep: 0x00000008)
uart_gcs_cnode = cnode (5 bits)
uart_gcs_fault_ep = ep
uart_gcs_group_bin_pd = pd
uart_gcs_interface_init_ep = ep
uart_gcs_post_init_ep = ep
uart_gcs_pre_init_ep = ep
uart_gcs_read_sem = ep
uart_gcs_write_sem = ep
uart_inf_ep = ep
uart_px4_8_0_control_9_tcb = tcb (addr: 0x13de00, ip: 0x159b0, sp: 0x156000, elf: uart_px4_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [3], fault_ep: 0x00000004)
uart_px4_8_0_fault_handler_15_0000_tcb = tcb (addr: 0x134e00, ip: 0x159b0, sp: 0x144000, elf: uart_px4_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [9])
uart_px4_8_interrupt_9_0000_tcb = tcb (addr: 0x13ae00, ip: 0x159b0, sp: 0x150000, elf: uart_px4_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [5], fault_ep: 0x00000006)
uart_px4_8_uart_4_0000_tcb = tcb (addr: 0x137e00, ip: 0x159b0, sp: 0x14a000, elf: uart_px4_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [7], fault_ep: 0x00000008)
uart_px4_cnode = cnode (5 bits)
uart_px4_fault_ep = ep
uart_px4_group_bin_pd = pd
uart_px4_interface_init_ep = ep
uart_px4_post_init_ep = ep
uart_px4_pre_init_ep = ep
uart_px4_read_sem = ep
uart_px4_write_sem = ep
uartbase_irq_irq = irq
uartbase_irq_ntfn = notification
uartpx4_inf_ep = ep
uartpx4_irq_irq = irq
uartpx4_irq_ntfn = notification
vm_2_0_control_9_tcb = tcb (addr: 0x5ae3e00, ip: 0x379fc, sp: 0x5af6000, elf: vm_group_bin, prio: 101,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [2], fault_ep: 0x00000003)
vm_2_0_fault_handler_15_0000_tcb = tcb (addr: 0x5adde00, ip: 0x379fc, sp: 0x5aea000, elf: vm_group_bin, prio: 255,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [6])
vm_2_restart_event_13_0000_tcb = tcb (addr: 0x5ae0e00, ip: 0x379fc, sp: 0x5af0000, elf: vm_group_bin, prio: 254,                max_prio: 254, crit: 1, max_crit: 1,                affinity: 0, init: [4], fault_ep: 0x00000005)
vm_asid_pool = asid_pool
vm_cnode = cnode (23 bits)
vm_fault_ep = ep
vm_group_bin_pd = pd
vm_interface_init_ep = ep
vm_irq_103 = irq
vm_irq_107 = irq
vm_irq_109 = irq
vm_irq_27 = irq
vm_irq_85 = irq
vm_irq_notification_obj = notification
vm_mmio_frame_268500992 = frame (4k, paddr: 0x10010000)
vm_mmio_frame_268517376 = frame (4k, paddr: 0x10014000)
vm_mmio_frame_268566528 = frame (4k, paddr: 0x10020000)
vm_mmio_frame_322961408 = frame (4k, paddr: 0x13400000)
vm_post_init_ep = ep
vm_pre_init_ep = ep
vm_simple_untyped_24_pool_0 = ut (24 bits)
vm_simple_untyped_24_pool_1 = ut (24 bits)
vm_simple_untyped_24_pool_2 = ut (24 bits)
vm_simple_untyped_24_pool_3 = ut (24 bits)
vm_simple_untyped_24_pool_4 = ut (24 bits)
vm_simple_untyped_24_pool_5 = ut (24 bits)
vm_simple_untyped_24_pool_6 = ut (24 bits)
vm_simple_untyped_24_pool_7 = ut (24 bits)
vm_simple_untyped_24_pool_8 = ut (24 bits)
vm_simple_untyped_24_pool_9 = ut (24 bits)
vm_untyped_cap_1073741824 = ut (29 bits, paddr: 0x40000000)
vm_untyped_cap_268435456 = ut (12 bits, paddr: 0x10000000)
vm_untyped_cap_268533760 = ut (12 bits, paddr: 0x10018000)
vm_untyped_cap_268550144 = ut (12 bits, paddr: 0x1001c000)
vm_untyped_cap_268632064 = ut (12 bits, paddr: 0x10030000)
vm_untyped_cap_268664832 = ut (12 bits, paddr: 0x10038000)
vm_untyped_cap_268697600 = ut (12 bits, paddr: 0x10040000)
vm_untyped_cap_268701696 = ut (12 bits, paddr: 0x10041000)
vm_untyped_cap_268705792 = ut (12 bits, paddr: 0x10042000)
vm_untyped_cap_268709888 = ut (12 bits, paddr: 0x10043000)
vm_untyped_cap_268713984 = ut (12 bits, paddr: 0x10044000)
vm_untyped_cap_268763136 = ut (12 bits, paddr: 0x10050000)
vm_untyped_cap_273178624 = ut (12 bits, paddr: 0x10486000)
vm_untyped_cap_303104000 = ut (12 bits, paddr: 0x12110000)
vm_untyped_cap_303235072 = ut (12 bits, paddr: 0x12130000)
vm_untyped_cap_304087040 = ut (12 bits, paddr: 0x12200000)
vm_untyped_cap_304218112 = ut (12 bits, paddr: 0x12220000)
vm_untyped_cap_314703872 = ut (12 bits, paddr: 0x12c20000)
vm_vm_sem = ep
}

caps {
can_obj_7_0_control_9_tcb {
cspace: can_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_can_obj_group_bin_0226 (RW)
vspace: can_obj_group_bin_pd
}
can_obj_7_0_fault_handler_15_0000_tcb {
cspace: can_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_can_obj_group_bin_0084 (RW)
vspace: can_obj_group_bin_pd
}
can_obj_7_Int_3_0000_tcb {
cspace: can_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_can_obj_group_bin_0085 (RW)
vspace: can_obj_group_bin_pd
}
can_obj_cnode {
0x1: can_obj_m_test (RW)
0x2: can_obj_7_0_control_9_tcb
0x3: can_obj_fault_ep (RWX, badge: 2)
0x4: can_obj_7_Int_3_0000_tcb
0x5: can_obj_fault_ep (RWX, badge: 4)
0x6: can_obj_7_0_fault_handler_15_0000_tcb
0x7: can_obj_fault_ep (RWX)
0x8: can_obj_pre_init_ep (RW)
0x9: can_obj_interface_init_ep (RW)
0xa: can_obj_post_init_ep (RW)
0xb: can_spi_ep (WX, badge: 0)
0xc: gpio_can_int_notification_0 (R)
0xd: gpio_can_int_handoff_0 (RW)
0xe: gpio_can_int_lock_0 (RW)
0xf: gpio_can_intAck_notification_0 (W)
}
can_obj_group_bin_pd {
0x0: pt_can_obj_group_bin_0000
}
clk_obj_7_0_control_9_tcb {
cspace: clk_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_clk_obj_group_bin_0227 (RW)
vspace: clk_obj_group_bin_pd
}
clk_obj_7_0_fault_handler_15_0000_tcb {
cspace: clk_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_clk_obj_group_bin_0084 (RW)
vspace: clk_obj_group_bin_pd
}
clk_obj_7_clktree_7_0000_tcb {
cspace: clk_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_clk_obj_group_bin_0085 (RW)
vspace: clk_obj_group_bin_pd
}
clk_obj_cnode {
0x1: clk_obj_7_0_control_9_tcb
0x2: clk_obj_fault_ep (RWX, badge: 1)
0x3: clk_obj_7_clktree_7_0000_tcb
0x4: clk_obj_fault_ep (RWX, badge: 3)
0x5: clk_obj_7_0_fault_handler_15_0000_tcb
0x6: clk_obj_fault_ep (RWX)
0x7: clk_obj_pre_init_ep (RW)
0x8: clk_obj_interface_init_ep (RW)
0x9: clk_obj_post_init_ep (RW)
0xa: spi_clk_ep (RW)
}
clk_obj_group_bin_pd {
0x0: pt_clk_obj_group_bin_0000
0x1: pt_clk_obj_group_bin_0106
0x2: pt_clk_obj_group_bin_0285
}
gpio_grp26_irq_irq {
0x0: gpio_grp26_irq_ntfn (R)
}
gpio_grp28_irq_irq {
0x0: gpio_grp28_irq_ntfn (R)
}
gpio_grp31_irq_irq {
0x0: gpio_grp31_irq_ntfn (R)
}
gpio_obj_8_0_control_9_tcb {
cspace: gpio_obj_cnode (guard: 0, guard_size: 26)
ipc_buffer_slot: frame_gpio_obj_group_bin_0260 (RW)
vspace: gpio_obj_group_bin_pd
}
gpio_obj_8_0_fault_handler_15_0000_tcb {
cspace: gpio_obj_cnode (guard: 0, guard_size: 26)
ipc_buffer_slot: frame_gpio_obj_group_bin_0042 (RW)
vspace: gpio_obj_group_bin_pd
}
gpio_obj_8_CANIntAck_9_0000_tcb {
cspace: gpio_obj_cnode (guard: 0, guard_size: 26)
ipc_buffer_slot: frame_gpio_obj_group_bin_0024 (RW)
vspace: gpio_obj_group_bin_pd
}
gpio_obj_8_gpio_4_0000_tcb {
cspace: gpio_obj_cnode (guard: 0, guard_size: 26)
ipc_buffer_slot: frame_gpio_obj_group_bin_0004 (RW)
vspace: gpio_obj_group_bin_pd
}
gpio_obj_8_irq_grp26_int_13_0000_tcb {
cspace: gpio_obj_cnode (guard: 0, guard_size: 26)
ipc_buffer_slot: frame_gpio_obj_group_bin_0297 (RW)
vspace: gpio_obj_group_bin_pd
}
gpio_obj_8_irq_grp28_int_13_0000_tcb {
cspace: gpio_obj_cnode (guard: 0, guard_size: 26)
ipc_buffer_slot: frame_gpio_obj_group_bin_0277 (RW)
vspace: gpio_obj_group_bin_pd
}
gpio_obj_8_irq_grp31_int_13_0000_tcb {
cspace: gpio_obj_cnode (guard: 0, guard_size: 26)
ipc_buffer_slot: frame_gpio_obj_group_bin_0318 (RW)
vspace: gpio_obj_group_bin_pd
}
gpio_obj_8_xint16_31_int_13_0000_tcb {
cspace: gpio_obj_cnode (guard: 0, guard_size: 26)
ipc_buffer_slot: frame_gpio_obj_group_bin_0339 (RW)
vspace: gpio_obj_group_bin_pd
}
gpio_obj_cnode {
0x10: gpio_obj_fault_ep (RWX)
0x11: gpio_obj_pre_init_ep (RW)
0x12: gpio_obj_interface_init_ep (RW)
0x13: gpio_obj_post_init_ep (RW)
0x14: gpio_grp28_irq_ntfn (R)
0x15: gpio_grp28_irq_irq
0x16: gpio_grp26_irq_ntfn (R)
0x17: gpio_grp26_irq_irq
0x18: gpio_grp31_irq_ntfn (R)
0x19: gpio_grp31_irq_irq
0x1: gpio_obj_8_0_control_9_tcb
0x1a: gpio_xint16_31_irq_ntfn (R)
0x1b: gpio_xint16_31_irq_irq
0x1c: spi_gpio_ep (RW)
0x1d: gpio_obj_cnode (guard: 0, guard_size: 26)
0x1f: gpio_can_int_notification_0 (W)
0x20: gpio_can_intAck_notification_0 (R)
0x21: gpio_can_intAck_handoff_0 (RW)
0x22: gpio_can_intAck_lock_0 (RW)
0x2: gpio_obj_fault_ep (RWX, badge: 1)
0x3: gpio_obj_8_irq_grp28_int_13_0000_tcb
0x4: gpio_obj_fault_ep (RWX, badge: 3)
0x5: gpio_obj_8_irq_grp26_int_13_0000_tcb
0x6: gpio_obj_fault_ep (RWX, badge: 5)
0x7: gpio_obj_8_irq_grp31_int_13_0000_tcb
0x8: gpio_obj_fault_ep (RWX, badge: 7)
0x9: gpio_obj_8_xint16_31_int_13_0000_tcb
0xa: gpio_obj_fault_ep (RWX, badge: 9)
0xb: gpio_obj_8_gpio_4_0000_tcb
0xc: gpio_obj_fault_ep (RWX, badge: 11)
0xd: gpio_obj_8_CANIntAck_9_0000_tcb
0xe: gpio_obj_fault_ep (RWX, badge: 13)
0xf: gpio_obj_8_0_fault_handler_15_0000_tcb
}
gpio_obj_group_bin_pd {
0x0: pt_gpio_obj_group_bin_0000
0x1: pt_gpio_obj_group_bin_0007
0x2: pt_gpio_obj_group_bin_0052
}
gpio_xint16_31_irq_irq {
0x0: gpio_xint16_31_irq_ntfn (R)
}
i2c0_irq_irq {
0x0: i2c0_irq_ntfn (R)
}
pilot_obj_9_0_control_9_tcb {
cspace: pilot_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pilot_obj_group_bin_0207 (RW)
vspace: pilot_obj_group_bin_pd
}
pilot_obj_9_0_fault_handler_15_0000_tcb {
cspace: pilot_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pilot_obj_group_bin_0260 (RW)
vspace: pilot_obj_group_bin_pd
}
pilot_obj_9_mavlink_7_0000_tcb {
cspace: pilot_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pilot_obj_group_bin_0096 (RW)
vspace: pilot_obj_group_bin_pd
}
pilot_obj_cnode {
0x11: fd_pwm.vm_pwm_ep (WX, badge: 0)
0x1: pilot_obj_9_0_control_9_tcb
0x2: pilot_obj_fault_ep (RWX, badge: 1)
0x3: pilot_obj_9_mavlink_7_0000_tcb
0x4: pilot_obj_fault_ep (RWX, badge: 3)
0x5: pilot_obj_9_0_fault_handler_15_0000_tcb
0x6: pilot_obj_fault_ep (RWX)
0x7: pilot_obj_pre_init_ep (RW)
0x8: pilot_obj_interface_init_ep (RW)
0x9: pilot_obj_post_init_ep (RW)
0xa: uart_inf_ep (WX, badge: 0)
0xb: uartpx4_inf_ep (WX, badge: 0)
0xc: pwm_sig_notification_0 (W)
0xd: restart_vm_notification_0 (W)
0xe: gcs_recv_inf.px4_recv_inf_ep (RW)
0xf: pilot_obj_cnode (guard: 0, guard_size: 27)
}
pilot_obj_group_bin_pd {
0x0: pt_pilot_obj_group_bin_0000
}
pt_can_obj_group_bin_0000 {
0x100: frame_can_obj_group_bin_0112 (RW)
0x101: frame_can_obj_group_bin_0202 (RW)
0x102: frame_can_obj_group_bin_0289 (RW)
0x103: frame_can_obj_group_bin_0072 (RW)
0x104: frame_can_obj_group_bin_0162 (RW)
0x105: frame_can_obj_group_bin_0249 (RW)
0x106: frame_can_obj_group_bin_0033 (RW)
0x107: frame_can_obj_group_bin_0119 (RW)
0x108: frame_can_obj_group_bin_0208 (RW)
0x109: frame_can_obj_group_bin_0295 (RW)
0x10: frame_can_obj_group_bin_0000 (RX)
0x10a: frame_can_obj_group_bin_0079 (RW)
0x10b: frame_can_obj_group_bin_0168 (RW)
0x10c: frame_can_obj_group_bin_0256 (RW)
0x10d: frame_can_obj_group_bin_0039 (RW)
0x10e: frame_can_obj_group_bin_0126 (RW)
0x10f: frame_can_obj_group_bin_0215 (RW)
0x110: frame_can_obj_group_bin_0302 (RW)
0x111: frame_can_obj_group_bin_0087 (RW)
0x112: frame_can_obj_group_bin_0174 (RW)
0x113: frame_can_obj_group_bin_0263 (RW)
0x114: frame_can_obj_group_bin_0046 (RW)
0x115: frame_can_obj_group_bin_0134 (RW)
0x116: frame_can_obj_group_bin_0223 (RW)
0x117: frame_can_obj_group_bin_0006 (RW)
0x118: frame_can_obj_group_bin_0171 (RW)
0x119: frame_can_obj_group_bin_0163 (RW)
0x11: frame_can_obj_group_bin_0001 (RX)
0x11a: frame_can_obj_group_bin_0073 (RW)
0x11b: frame_can_obj_group_bin_0273 (RW)
0x11c: frame_can_obj_group_bin_0103 (RW)
0x11d: frame_can_obj_group_bin_0241 (RW)
0x11e: frame_can_obj_group_bin_0070 (RW)
0x11f: frame_can_obj_group_bin_0206 (RW)
0x120: frame_can_obj_group_bin_0040 (RW)
0x121: frame_can_obj_group_bin_0060 (RW)
0x122: frame_can_obj_group_bin_0153 (RW)
0x123: frame_can_obj_group_bin_0142 (RW)
0x124: frame_can_obj_group_bin_0240 (RW)
0x125: frame_can_obj_group_bin_0108 (RW)
0x126: frame_can_obj_group_bin_0012 (RW)
0x127: frame_can_obj_group_bin_0051 (RW)
0x128: frame_can_obj_group_bin_0287 (RW)
0x129: frame_can_obj_group_bin_0225 (RW)
0x12: frame_can_obj_group_bin_0214 (RX)
0x12a: frame_can_obj_group_bin_0160 (RW)
0x12b: frame_can_obj_group_bin_0247 (RW)
0x12c: frame_can_obj_group_bin_0031 (RW)
0x12d: frame_can_obj_group_bin_0117 (RW)
0x12e: frame_can_obj_group_bin_0211 (RW)
0x12f: frame_can_obj_group_bin_0293 (RW)
0x130: frame_can_obj_group_bin_0077 (RW)
0x131: frame_can_obj_group_bin_0183 (RW)
0x132: frame_can_obj_group_bin_0252 (RW)
0x134: frame_can_obj_group_bin_0084 (RW)
0x137: frame_can_obj_group_bin_0085 (RW)
0x13: frame_can_obj_group_bin_0292 (RX)
0x13a: frame_can_obj_group_bin_0226 (RW)
0x13d: frame_can_obj_group_bin_0025 (RW)
0x13e: frame_can_obj_group_bin_0180 (RW)
0x13f: frame_can_obj_group_bin_0250 (RW)
0x140: frame_can_obj_group_bin_0270 (RW)
0x143: frame_can_obj_group_bin_0231 (RW)
0x144: frame_can_obj_group_bin_0015 (RW)
0x145: frame_can_obj_group_bin_0100 (RW)
0x146: frame_can_obj_group_bin_0191 (RW)
0x149: frame_can_obj_group_bin_0149 (RW)
0x14: frame_can_obj_group_bin_0067 (RX)
0x14a: frame_can_obj_group_bin_0123 (RW)
0x14b: frame_can_obj_group_bin_0022 (RW)
0x14c: frame_can_obj_group_bin_0107 (RW)
0x14e: frame_can_obj_group_bin_0284 (RWX)
0x15: frame_can_obj_group_bin_0146 (RX)
0x16: frame_can_obj_group_bin_0224 (RX)
0x17: frame_can_obj_group_bin_0300 (RX)
0x18: frame_can_obj_group_bin_0076 (RX)
0x19: frame_can_obj_group_bin_0080 (RX)
0x1a: frame_can_obj_group_bin_0157 (RX)
0x1b: frame_can_obj_group_bin_0007 (RX)
0x1c: frame_can_obj_group_bin_0086 (RX)
0x1d: frame_can_obj_group_bin_0165 (RX)
0x1e: frame_can_obj_group_bin_0243 (RX)
0x1f: frame_can_obj_group_bin_0018 (RX)
0x20: frame_can_obj_group_bin_0094 (RX)
0x30: frame_can_obj_group_bin_0004 (RW)
0x31: frame_can_obj_group_bin_0212 (RW)
0x32: frame_can_obj_group_bin_0290 (RW)
0x33: frame_can_obj_group_bin_0065 (RW)
0x34: frame_can_obj_group_bin_0143 (RW)
0x35: frame_can_obj_group_bin_0221 (RW)
0x36: frame_can_obj_group_bin_0298 (RW)
0x37: frame_can_obj_group_bin_0074 (RW)
0x38: frame_can_obj_group_bin_0152 (RW)
0x39: frame_can_obj_group_bin_0232 (RW)
0x3a: frame_can_obj_group_bin_0005 (RW)
0x3b: frame_can_obj_group_bin_0083 (RW)
0x3c: frame_can_obj_group_bin_0164 (RW)
0x3d: frame_can_obj_group_bin_0242 (RW)
0x3e: frame_can_obj_group_bin_0016 (RW)
0x3f: frame_can_obj_group_bin_0092 (RW)
0x40: frame_can_obj_group_bin_0172 (RW)
0x41: frame_can_obj_group_bin_0251 (RW)
0x42: frame_can_obj_group_bin_0026 (RW)
0x43: frame_can_obj_group_bin_0102 (RW)
0x44: frame_can_obj_group_bin_0181 (RW)
0x45: frame_can_obj_group_bin_0260 (RW)
0x46: frame_can_obj_group_bin_0034 (RW)
0x47: frame_can_obj_group_bin_0111 (RW)
0x48: frame_can_obj_group_bin_0192 (RW)
0x49: frame_can_obj_group_bin_0269 (RW)
0x4a: frame_can_obj_group_bin_0043 (RW)
0x4b: frame_can_obj_group_bin_0120 (RW)
0x4c: frame_can_obj_group_bin_0201 (RW)
0x4d: frame_can_obj_group_bin_0279 (RW)
0x4e: frame_can_obj_group_bin_0053 (RW)
0x4f: frame_can_obj_group_bin_0130 (RW)
0x50: frame_can_obj_group_bin_0209 (RW)
0x51: frame_can_obj_group_bin_0288 (RW)
0x52: frame_can_obj_group_bin_0063 (RW)
0x53: frame_can_obj_group_bin_0140 (RW)
0x54: frame_can_obj_group_bin_0219 (RW)
0x55: frame_can_obj_group_bin_0296 (RW)
0x56: frame_can_obj_group_bin_0071 (RW)
0x57: frame_can_obj_group_bin_0150 (RW)
0x58: frame_can_obj_group_bin_0230 (RW)
0x59: frame_can_obj_group_bin_0002 (RW)
0x5a: frame_can_obj_group_bin_0081 (RW)
0x5b: frame_can_obj_group_bin_0161 (RW)
0x5c: frame_can_obj_group_bin_0239 (RW)
0x5d: frame_can_obj_group_bin_0014 (RW)
0x5e: frame_can_obj_group_bin_0090 (RW)
0x5f: frame_can_obj_group_bin_0169 (RW)
0x60: frame_can_obj_group_bin_0248 (RW)
0x61: frame_can_obj_group_bin_0023 (RW)
0x62: frame_can_obj_group_bin_0099 (RW)
0x63: frame_can_obj_group_bin_0178 (RW)
0x64: frame_can_obj_group_bin_0257 (RW)
0x65: frame_can_obj_group_bin_0032 (RW)
0x66: frame_can_obj_group_bin_0109 (RW)
0x67: frame_can_obj_group_bin_0234 (RW)
0x68: frame_can_obj_group_bin_0267 (RW)
0x69: frame_can_obj_group_bin_0041 (RW)
0x6a: frame_can_obj_group_bin_0118 (RW)
0x6b: frame_can_obj_group_bin_0199 (RW)
0x6c: frame_can_obj_group_bin_0277 (RW)
0x6d: frame_can_obj_group_bin_0050 (RW)
0x6e: frame_can_obj_group_bin_0127 (RW)
0x6f: frame_can_obj_group_bin_0207 (RW)
0x70: frame_can_obj_group_bin_0285 (RW)
0x71: frame_can_obj_group_bin_0061 (RW)
0x72: frame_can_obj_group_bin_0137 (RW)
0x73: frame_can_obj_group_bin_0216 (RW)
0x74: frame_can_obj_group_bin_0294 (RW)
0x75: frame_can_obj_group_bin_0069 (RW)
0x76: frame_can_obj_group_bin_0148 (RW)
0x77: frame_can_obj_group_bin_0228 (RW)
0x78: frame_can_obj_group_bin_0303 (RW)
0x79: frame_can_obj_group_bin_0078 (RW)
0x7a: frame_can_obj_group_bin_0158 (RW)
0x7b: frame_can_obj_group_bin_0237 (RW)
0x7c: frame_can_obj_group_bin_0011 (RW)
0x7d: frame_can_obj_group_bin_0088 (RW)
0x7e: frame_can_obj_group_bin_0167 (RW)
0x7f: frame_can_obj_group_bin_0245 (RW)
0x80: frame_can_obj_group_bin_0021 (RW)
0x81: frame_can_obj_group_bin_0097 (RW)
0x82: frame_can_obj_group_bin_0175 (RW)
0x83: frame_can_obj_group_bin_0255 (RW)
0x84: frame_can_obj_group_bin_0029 (RW)
0x85: frame_can_obj_group_bin_0106 (RW)
0x86: frame_can_obj_group_bin_0187 (RW)
0x87: frame_can_obj_group_bin_0264 (RW)
0x88: frame_can_obj_group_bin_0038 (RW)
0x89: frame_can_obj_group_bin_0115 (RW)
0x8a: frame_can_obj_group_bin_0197 (RW)
0x8b: frame_can_obj_group_bin_0275 (RW)
0x8c: frame_can_obj_group_bin_0047 (RW)
0x8d: frame_can_obj_group_bin_0125 (RW)
0x8e: frame_can_obj_group_bin_0205 (RW)
0x8f: frame_can_obj_group_bin_0283 (RW)
0x90: frame_can_obj_group_bin_0058 (RW)
0x91: frame_can_obj_group_bin_0135 (RW)
0x92: frame_can_obj_group_bin_0166 (RW)
0x93: frame_can_obj_group_bin_0254 (RW)
0x94: frame_can_obj_group_bin_0037 (RW)
0x95: frame_can_obj_group_bin_0124 (RW)
0x96: frame_can_obj_group_bin_0213 (RW)
0x97: frame_can_obj_group_bin_0299 (RW)
0x98: frame_can_obj_group_bin_0121 (RW)
0x99: frame_can_obj_group_bin_0156 (RW)
0x9a: frame_can_obj_group_bin_0235 (RW)
0x9b: frame_can_obj_group_bin_0045 (RW)
0x9c: frame_can_obj_group_bin_0132 (RW)
0x9d: frame_can_obj_group_bin_0193 (RW)
0x9e: frame_can_obj_group_bin_0024 (RW)
0x9f: frame_can_obj_group_bin_0159 (RW)
0xa0: frame_can_obj_group_bin_0182 (RW)
0xa1: frame_can_obj_group_bin_0173 (RW)
0xa2: frame_can_obj_group_bin_0253 (RW)
0xa3: frame_can_obj_group_bin_0027 (RW)
0xa4: frame_can_obj_group_bin_0104 (RW)
0xa5: frame_can_obj_group_bin_0184 (RW)
0xa6: frame_can_obj_group_bin_0262 (RW)
0xa7: frame_can_obj_group_bin_0036 (RW)
0xa8: frame_can_obj_group_bin_0113 (RW)
0xa9: frame_can_obj_group_bin_0195 (RW)
0xaa: frame_can_obj_group_bin_0272 (RW)
0xab: frame_can_obj_group_bin_0238 (RW)
0xac: frame_can_obj_group_bin_0122 (RW)
0xad: frame_can_obj_group_bin_0203 (RW)
0xae: frame_can_obj_group_bin_0281 (RW)
0xaf: frame_can_obj_group_bin_0055 (RW)
0xb0: frame_can_obj_group_bin_0068 (RW)
0xb1: frame_can_obj_group_bin_0246 (RW)
0xb2: frame_can_obj_group_bin_0244 (RW)
0xb3: frame_can_obj_group_bin_0028 (RW)
0xb4: frame_can_obj_group_bin_0114 (RW)
0xb5: frame_can_obj_group_bin_0204 (RW)
0xb6: frame_can_obj_group_bin_0291 (RW)
0xb7: frame_can_obj_group_bin_0075 (RW)
0xb8: frame_can_obj_group_bin_0210 (RW)
0xb9: frame_can_obj_group_bin_0042 (RW)
0xba: frame_can_obj_group_bin_0176 (RW)
0xbb: frame_can_obj_group_bin_0008 (RW)
0xbc: frame_can_obj_group_bin_0144 (RW)
0xbd: frame_can_obj_group_bin_0280 (RW)
0xbe: frame_can_obj_group_bin_0110 (RW)
0xbf: frame_can_obj_group_bin_0009 (RW)
0xc0: frame_can_obj_group_bin_0261 (RW)
0xc1: frame_can_obj_group_bin_0044 (RW)
0xc2: frame_can_obj_group_bin_0131 (RW)
0xc3: frame_can_obj_group_bin_0220 (RW)
0xc4: frame_can_obj_group_bin_0003 (RW)
0xc5: frame_can_obj_group_bin_0091 (RW)
0xc6: frame_can_obj_group_bin_0179 (RW)
0xc7: frame_can_obj_group_bin_0268 (RW)
0xc8: frame_can_obj_group_bin_0052 (RW)
0xc9: frame_can_obj_group_bin_0138 (RW)
0xca: frame_can_obj_group_bin_0229 (RW)
0xcb: frame_can_obj_group_bin_0013 (RW)
0xcc: frame_can_obj_group_bin_0098 (RW)
0xcd: frame_can_obj_group_bin_0189 (RW)
0xce: frame_can_obj_group_bin_0276 (RW)
0xcf: frame_can_obj_group_bin_0059 (RW)
0xd0: frame_can_obj_group_bin_0147 (RW)
0xd1: frame_can_obj_group_bin_0236 (RW)
0xd2: frame_can_obj_group_bin_0020 (RW)
0xd3: frame_can_obj_group_bin_0105 (RW)
0xd4: frame_can_obj_group_bin_0196 (RW)
0xd5: frame_can_obj_group_bin_0282 (RW)
0xd6: frame_can_obj_group_bin_0066 (RW)
0xd7: frame_can_obj_group_bin_0155 (RW)
0xd8: frame_can_obj_group_bin_0297 (RW)
0xd9: frame_can_obj_group_bin_0128 (RW)
0xda: frame_can_obj_group_bin_0265 (RW)
0xdb: frame_can_obj_group_bin_0095 (RW)
0xdc: frame_can_obj_group_bin_0233 (RW)
0xdd: frame_can_obj_group_bin_0064 (RW)
0xde: frame_can_obj_group_bin_0200 (RW)
0xdf: frame_can_obj_group_bin_0030 (RW)
0xe0: frame_can_obj_group_bin_0035 (RW)
0xe1: frame_can_obj_group_bin_0301 (RW)
0xe2: frame_can_obj_group_bin_0133 (RW)
0xe3: frame_can_obj_group_bin_0271 (RW)
0xe4: frame_can_obj_group_bin_0082 (RW)
0xe5: frame_can_obj_group_bin_0170 (RW)
0xe6: frame_can_obj_group_bin_0258 (RW)
0xe7: frame_can_obj_group_bin_0190 (RW)
0xe8: frame_can_obj_group_bin_0129 (RW)
0xe9: frame_can_obj_group_bin_0218 (RW)
0xea: frame_can_obj_group_bin_0093 (RW)
0xeb: frame_can_obj_group_bin_0089 (RW)
0xec: frame_can_obj_group_bin_0177 (RW)
0xed: frame_can_obj_group_bin_0266 (RW)
0xee: frame_can_obj_group_bin_0049 (RW)
0xef: frame_can_obj_group_bin_0136 (RW)
0xf0: frame_can_obj_group_bin_0227 (RW)
0xf1: frame_can_obj_group_bin_0010 (RW)
0xf2: frame_can_obj_group_bin_0096 (RW)
0xf3: frame_can_obj_group_bin_0186 (RW)
0xf4: frame_can_obj_group_bin_0274 (RW)
0xf5: frame_can_obj_group_bin_0057 (RW)
0xf6: frame_can_obj_group_bin_0145 (RW)
0xf7: frame_can_obj_group_bin_0019 (RW)
0xf8: frame_can_obj_group_bin_0101 (RW)
0xf9: frame_can_obj_group_bin_0217 (RW)
0xfa: frame_can_obj_group_bin_0048 (RW)
0xfb: frame_can_obj_group_bin_0185 (RW)
0xfc: frame_can_obj_group_bin_0017 (RW)
0xfd: frame_can_obj_group_bin_0151 (RW)
0xfe: frame_can_obj_group_bin_0286 (RW)
0xff: frame_can_obj_group_bin_0116 (RW)
}
pt_clk_obj_group_bin_0000 {
0x100: frame_clk_obj_group_bin_0113 (RW)
0x101: frame_clk_obj_group_bin_0203 (RW)
0x102: frame_clk_obj_group_bin_0291 (RW)
0x103: frame_clk_obj_group_bin_0072 (RW)
0x104: frame_clk_obj_group_bin_0163 (RW)
0x105: frame_clk_obj_group_bin_0251 (RW)
0x106: frame_clk_obj_group_bin_0033 (RW)
0x107: frame_clk_obj_group_bin_0120 (RW)
0x108: frame_clk_obj_group_bin_0209 (RW)
0x109: frame_clk_obj_group_bin_0297 (RW)
0x10: frame_clk_obj_group_bin_0000 (RX)
0x10a: frame_clk_obj_group_bin_0079 (RW)
0x10b: frame_clk_obj_group_bin_0169 (RW)
0x10c: frame_clk_obj_group_bin_0258 (RW)
0x10d: frame_clk_obj_group_bin_0039 (RW)
0x10e: frame_clk_obj_group_bin_0127 (RW)
0x10f: frame_clk_obj_group_bin_0216 (RW)
0x110: frame_clk_obj_group_bin_0304 (RW)
0x111: frame_clk_obj_group_bin_0087 (RW)
0x112: frame_clk_obj_group_bin_0175 (RW)
0x113: frame_clk_obj_group_bin_0265 (RW)
0x114: frame_clk_obj_group_bin_0046 (RW)
0x115: frame_clk_obj_group_bin_0135 (RW)
0x116: frame_clk_obj_group_bin_0224 (RW)
0x117: frame_clk_obj_group_bin_0006 (RW)
0x118: frame_clk_obj_group_bin_0172 (RW)
0x119: frame_clk_obj_group_bin_0164 (RW)
0x11: frame_clk_obj_group_bin_0001 (RX)
0x11a: frame_clk_obj_group_bin_0073 (RW)
0x11b: frame_clk_obj_group_bin_0275 (RW)
0x11c: frame_clk_obj_group_bin_0103 (RW)
0x11d: frame_clk_obj_group_bin_0243 (RW)
0x11e: frame_clk_obj_group_bin_0070 (RW)
0x11f: frame_clk_obj_group_bin_0207 (RW)
0x120: frame_clk_obj_group_bin_0040 (RW)
0x121: frame_clk_obj_group_bin_0060 (RW)
0x122: frame_clk_obj_group_bin_0154 (RW)
0x123: frame_clk_obj_group_bin_0143 (RW)
0x124: frame_clk_obj_group_bin_0242 (RW)
0x125: frame_clk_obj_group_bin_0109 (RW)
0x126: frame_clk_obj_group_bin_0012 (RW)
0x127: frame_clk_obj_group_bin_0051 (RW)
0x128: frame_clk_obj_group_bin_0289 (RW)
0x129: frame_clk_obj_group_bin_0226 (RW)
0x12: frame_clk_obj_group_bin_0215 (RX)
0x12a: frame_clk_obj_group_bin_0161 (RW)
0x12b: frame_clk_obj_group_bin_0249 (RW)
0x12c: frame_clk_obj_group_bin_0031 (RW)
0x12d: frame_clk_obj_group_bin_0118 (RW)
0x12e: frame_clk_obj_group_bin_0212 (RW)
0x12f: frame_clk_obj_group_bin_0295 (RW)
0x130: frame_clk_obj_group_bin_0077 (RW)
0x131: frame_clk_obj_group_bin_0184 (RW)
0x132: frame_clk_obj_group_bin_0254 (RW)
0x134: frame_clk_obj_group_bin_0084 (RW)
0x137: frame_clk_obj_group_bin_0085 (RW)
0x13: frame_clk_obj_group_bin_0294 (RX)
0x13a: frame_clk_obj_group_bin_0227 (RW)
0x13d: frame_clk_obj_group_bin_0025 (RW)
0x13e: frame_clk_obj_group_bin_0181 (RW)
0x13f: frame_clk_obj_group_bin_0252 (RW)
0x140: frame_clk_obj_group_bin_0272 (RW)
0x143: frame_clk_obj_group_bin_0232 (RW)
0x144: frame_clk_obj_group_bin_0015 (RW)
0x145: frame_clk_obj_group_bin_0100 (RW)
0x146: frame_clk_obj_group_bin_0192 (RW)
0x149: frame_clk_obj_group_bin_0150 (RW)
0x14: frame_clk_obj_group_bin_0067 (RX)
0x14a: frame_clk_obj_group_bin_0124 (RW)
0x14b: frame_clk_obj_group_bin_0022 (RW)
0x14c: frame_clk_obj_group_bin_0108 (RW)
0x15: frame_clk_obj_group_bin_0147 (RX)
0x16: frame_clk_obj_group_bin_0225 (RX)
0x17: frame_clk_obj_group_bin_0302 (RX)
0x18: frame_clk_obj_group_bin_0076 (RX)
0x19: frame_clk_obj_group_bin_0080 (RX)
0x1a: frame_clk_obj_group_bin_0158 (RX)
0x1b: frame_clk_obj_group_bin_0007 (RX)
0x1c: frame_clk_obj_group_bin_0086 (RX)
0x1d: frame_clk_obj_group_bin_0166 (RX)
0x1e: frame_clk_obj_group_bin_0245 (RX)
0x1f: frame_clk_obj_group_bin_0018 (RX)
0x20: frame_clk_obj_group_bin_0094 (RX)
0x30: frame_clk_obj_group_bin_0004 (RW)
0x31: frame_clk_obj_group_bin_0213 (RW)
0x32: frame_clk_obj_group_bin_0292 (RW)
0x33: frame_clk_obj_group_bin_0065 (RW)
0x34: frame_clk_obj_group_bin_0144 (RW)
0x35: frame_clk_obj_group_bin_0222 (RW)
0x36: frame_clk_obj_group_bin_0300 (RW)
0x37: frame_clk_obj_group_bin_0074 (RW)
0x38: frame_clk_obj_group_bin_0153 (RW)
0x39: frame_clk_obj_group_bin_0233 (RW)
0x3a: frame_clk_obj_group_bin_0005 (RW)
0x3b: frame_clk_obj_group_bin_0083 (RW)
0x3c: frame_clk_obj_group_bin_0165 (RW)
0x3d: frame_clk_obj_group_bin_0244 (RW)
0x3e: frame_clk_obj_group_bin_0016 (RW)
0x3f: frame_clk_obj_group_bin_0092 (RW)
0x40: frame_clk_obj_group_bin_0173 (RW)
0x41: frame_clk_obj_group_bin_0253 (RW)
0x42: frame_clk_obj_group_bin_0026 (RW)
0x43: frame_clk_obj_group_bin_0102 (RW)
0x44: frame_clk_obj_group_bin_0182 (RW)
0x45: frame_clk_obj_group_bin_0262 (RW)
0x46: frame_clk_obj_group_bin_0034 (RW)
0x47: frame_clk_obj_group_bin_0112 (RW)
0x48: frame_clk_obj_group_bin_0193 (RW)
0x49: frame_clk_obj_group_bin_0271 (RW)
0x4a: frame_clk_obj_group_bin_0043 (RW)
0x4b: frame_clk_obj_group_bin_0121 (RW)
0x4c: frame_clk_obj_group_bin_0202 (RW)
0x4d: frame_clk_obj_group_bin_0281 (RW)
0x4e: frame_clk_obj_group_bin_0053 (RW)
0x4f: frame_clk_obj_group_bin_0131 (RW)
0x50: frame_clk_obj_group_bin_0210 (RW)
0x51: frame_clk_obj_group_bin_0290 (RW)
0x52: frame_clk_obj_group_bin_0063 (RW)
0x53: frame_clk_obj_group_bin_0141 (RW)
0x54: frame_clk_obj_group_bin_0220 (RW)
0x55: frame_clk_obj_group_bin_0298 (RW)
0x56: frame_clk_obj_group_bin_0071 (RW)
0x57: frame_clk_obj_group_bin_0151 (RW)
0x58: frame_clk_obj_group_bin_0231 (RW)
0x59: frame_clk_obj_group_bin_0002 (RW)
0x5a: frame_clk_obj_group_bin_0081 (RW)
0x5b: frame_clk_obj_group_bin_0162 (RW)
0x5c: frame_clk_obj_group_bin_0241 (RW)
0x5d: frame_clk_obj_group_bin_0014 (RW)
0x5e: frame_clk_obj_group_bin_0090 (RW)
0x5f: frame_clk_obj_group_bin_0170 (RW)
0x60: frame_clk_obj_group_bin_0250 (RW)
0x61: frame_clk_obj_group_bin_0023 (RW)
0x62: frame_clk_obj_group_bin_0099 (RW)
0x63: frame_clk_obj_group_bin_0179 (RW)
0x64: frame_clk_obj_group_bin_0259 (RW)
0x65: frame_clk_obj_group_bin_0032 (RW)
0x66: frame_clk_obj_group_bin_0110 (RW)
0x67: frame_clk_obj_group_bin_0235 (RW)
0x68: frame_clk_obj_group_bin_0269 (RW)
0x69: frame_clk_obj_group_bin_0041 (RW)
0x6a: frame_clk_obj_group_bin_0119 (RW)
0x6b: frame_clk_obj_group_bin_0200 (RW)
0x6c: frame_clk_obj_group_bin_0279 (RW)
0x6d: frame_clk_obj_group_bin_0050 (RW)
0x6e: frame_clk_obj_group_bin_0128 (RW)
0x6f: frame_clk_obj_group_bin_0208 (RW)
0x70: frame_clk_obj_group_bin_0287 (RW)
0x71: frame_clk_obj_group_bin_0061 (RW)
0x72: frame_clk_obj_group_bin_0138 (RW)
0x73: frame_clk_obj_group_bin_0217 (RW)
0x74: frame_clk_obj_group_bin_0296 (RW)
0x75: frame_clk_obj_group_bin_0069 (RW)
0x76: frame_clk_obj_group_bin_0149 (RW)
0x77: frame_clk_obj_group_bin_0229 (RW)
0x78: frame_clk_obj_group_bin_0305 (RW)
0x79: frame_clk_obj_group_bin_0078 (RW)
0x7a: frame_clk_obj_group_bin_0159 (RW)
0x7b: frame_clk_obj_group_bin_0238 (RW)
0x7c: frame_clk_obj_group_bin_0011 (RW)
0x7d: frame_clk_obj_group_bin_0088 (RW)
0x7e: frame_clk_obj_group_bin_0168 (RW)
0x7f: frame_clk_obj_group_bin_0247 (RW)
0x80: frame_clk_obj_group_bin_0021 (RW)
0x81: frame_clk_obj_group_bin_0097 (RW)
0x82: frame_clk_obj_group_bin_0176 (RW)
0x83: frame_clk_obj_group_bin_0257 (RW)
0x84: frame_clk_obj_group_bin_0029 (RW)
0x85: frame_clk_obj_group_bin_0107 (RW)
0x86: frame_clk_obj_group_bin_0188 (RW)
0x87: frame_clk_obj_group_bin_0266 (RW)
0x88: frame_clk_obj_group_bin_0038 (RW)
0x89: frame_clk_obj_group_bin_0116 (RW)
0x8a: frame_clk_obj_group_bin_0198 (RW)
0x8b: frame_clk_obj_group_bin_0277 (RW)
0x8c: frame_clk_obj_group_bin_0047 (RW)
0x8d: frame_clk_obj_group_bin_0126 (RW)
0x8e: frame_clk_obj_group_bin_0206 (RW)
0x8f: frame_clk_obj_group_bin_0286 (RW)
0x90: frame_clk_obj_group_bin_0058 (RW)
0x91: frame_clk_obj_group_bin_0136 (RW)
0x92: frame_clk_obj_group_bin_0167 (RW)
0x93: frame_clk_obj_group_bin_0256 (RW)
0x94: frame_clk_obj_group_bin_0037 (RW)
0x95: frame_clk_obj_group_bin_0125 (RW)
0x96: frame_clk_obj_group_bin_0214 (RW)
0x97: frame_clk_obj_group_bin_0301 (RW)
0x98: frame_clk_obj_group_bin_0122 (RW)
0x99: frame_clk_obj_group_bin_0157 (RW)
0x9a: frame_clk_obj_group_bin_0236 (RW)
0x9b: frame_clk_obj_group_bin_0045 (RW)
0x9c: frame_clk_obj_group_bin_0133 (RW)
0x9d: frame_clk_obj_group_bin_0194 (RW)
0x9e: frame_clk_obj_group_bin_0024 (RW)
0x9f: frame_clk_obj_group_bin_0160 (RW)
0xa0: frame_clk_obj_group_bin_0183 (RW)
0xa1: frame_clk_obj_group_bin_0174 (RW)
0xa2: frame_clk_obj_group_bin_0255 (RW)
0xa3: frame_clk_obj_group_bin_0027 (RW)
0xa4: frame_clk_obj_group_bin_0104 (RW)
0xa5: frame_clk_obj_group_bin_0185 (RW)
0xa6: frame_clk_obj_group_bin_0264 (RW)
0xa7: frame_clk_obj_group_bin_0036 (RW)
0xa8: frame_clk_obj_group_bin_0114 (RW)
0xa9: frame_clk_obj_group_bin_0196 (RW)
0xaa: frame_clk_obj_group_bin_0274 (RW)
0xab: frame_clk_obj_group_bin_0240 (RW)
0xac: frame_clk_obj_group_bin_0123 (RW)
0xad: frame_clk_obj_group_bin_0204 (RW)
0xae: frame_clk_obj_group_bin_0284 (RW)
0xaf: frame_clk_obj_group_bin_0055 (RW)
0xb0: frame_clk_obj_group_bin_0068 (RW)
0xb1: frame_clk_obj_group_bin_0248 (RW)
0xb2: frame_clk_obj_group_bin_0246 (RW)
0xb3: frame_clk_obj_group_bin_0028 (RW)
0xb4: frame_clk_obj_group_bin_0115 (RW)
0xb5: frame_clk_obj_group_bin_0205 (RW)
0xb6: frame_clk_obj_group_bin_0293 (RW)
0xb7: frame_clk_obj_group_bin_0075 (RW)
0xb8: frame_clk_obj_group_bin_0211 (RW)
0xb9: frame_clk_obj_group_bin_0042 (RW)
0xba: frame_clk_obj_group_bin_0177 (RW)
0xbb: frame_clk_obj_group_bin_0008 (RW)
0xbc: frame_clk_obj_group_bin_0145 (RW)
0xbd: frame_clk_obj_group_bin_0282 (RW)
0xbe: frame_clk_obj_group_bin_0111 (RW)
0xbf: frame_clk_obj_group_bin_0009 (RW)
0xc0: frame_clk_obj_group_bin_0263 (RW)
0xc1: frame_clk_obj_group_bin_0044 (RW)
0xc2: frame_clk_obj_group_bin_0132 (RW)
0xc3: frame_clk_obj_group_bin_0221 (RW)
0xc4: frame_clk_obj_group_bin_0003 (RW)
0xc5: frame_clk_obj_group_bin_0091 (RW)
0xc6: frame_clk_obj_group_bin_0180 (RW)
0xc7: frame_clk_obj_group_bin_0270 (RW)
0xc8: frame_clk_obj_group_bin_0052 (RW)
0xc9: frame_clk_obj_group_bin_0139 (RW)
0xca: frame_clk_obj_group_bin_0230 (RW)
0xcb: frame_clk_obj_group_bin_0013 (RW)
0xcc: frame_clk_obj_group_bin_0098 (RW)
0xcd: frame_clk_obj_group_bin_0190 (RW)
0xce: frame_clk_obj_group_bin_0278 (RW)
0xcf: frame_clk_obj_group_bin_0059 (RW)
0xd0: frame_clk_obj_group_bin_0148 (RW)
0xd1: frame_clk_obj_group_bin_0237 (RW)
0xd2: frame_clk_obj_group_bin_0020 (RW)
0xd3: frame_clk_obj_group_bin_0106 (RW)
0xd4: frame_clk_obj_group_bin_0197 (RW)
0xd5: frame_clk_obj_group_bin_0285 (RW)
0xd6: frame_clk_obj_group_bin_0066 (RW)
0xd7: frame_clk_obj_group_bin_0156 (RW)
0xd8: frame_clk_obj_group_bin_0299 (RW)
0xd9: frame_clk_obj_group_bin_0129 (RW)
0xda: frame_clk_obj_group_bin_0267 (RW)
0xdb: frame_clk_obj_group_bin_0095 (RW)
0xdc: frame_clk_obj_group_bin_0234 (RW)
0xdd: frame_clk_obj_group_bin_0064 (RW)
0xde: frame_clk_obj_group_bin_0201 (RW)
0xdf: frame_clk_obj_group_bin_0030 (RW)
0xe0: frame_clk_obj_group_bin_0035 (RW)
0xe1: frame_clk_obj_group_bin_0303 (RW)
0xe2: frame_clk_obj_group_bin_0134 (RW)
0xe3: frame_clk_obj_group_bin_0273 (RW)
0xe4: frame_clk_obj_group_bin_0082 (RW)
0xe5: frame_clk_obj_group_bin_0171 (RW)
0xe6: frame_clk_obj_group_bin_0260 (RW)
0xe7: frame_clk_obj_group_bin_0191 (RW)
0xe8: frame_clk_obj_group_bin_0130 (RW)
0xe9: frame_clk_obj_group_bin_0219 (RW)
0xea: frame_clk_obj_group_bin_0093 (RW)
0xeb: frame_clk_obj_group_bin_0089 (RW)
0xec: frame_clk_obj_group_bin_0178 (RW)
0xed: frame_clk_obj_group_bin_0268 (RW)
0xee: frame_clk_obj_group_bin_0049 (RW)
0xef: frame_clk_obj_group_bin_0137 (RW)
0xf0: frame_clk_obj_group_bin_0228 (RW)
0xf1: frame_clk_obj_group_bin_0010 (RW)
0xf2: frame_clk_obj_group_bin_0096 (RW)
0xf3: frame_clk_obj_group_bin_0187 (RW)
0xf4: frame_clk_obj_group_bin_0276 (RW)
0xf5: frame_clk_obj_group_bin_0057 (RW)
0xf6: frame_clk_obj_group_bin_0146 (RW)
0xf7: frame_clk_obj_group_bin_0019 (RW)
0xf8: frame_clk_obj_group_bin_0101 (RW)
0xf9: frame_clk_obj_group_bin_0218 (RW)
0xfa: frame_clk_obj_group_bin_0048 (RW)
0xfb: frame_clk_obj_group_bin_0186 (RW)
0xfc: frame_clk_obj_group_bin_0017 (RW)
0xfd: frame_clk_obj_group_bin_0152 (RW)
0xfe: frame_clk_obj_group_bin_0288 (RW)
0xff: frame_clk_obj_group_bin_0117 (RW)
}
pt_clk_obj_group_bin_0106 {
0x0: frame_clk_obj_group_bin_0239 (RW, uncached)
0x100: frame_clk_obj_group_bin_0105 (RW, uncached)
}
pt_clk_obj_group_bin_0285 {
0x0: frame_clk_obj_group_bin_0283 (RW, uncached)
}
pt_gpio_obj_group_bin_0000 {
0x100: frame_gpio_obj_group_bin_0183 (RW)
0x101: frame_gpio_obj_group_bin_0293 (RW)
0x102: frame_gpio_obj_group_bin_0052 (RW)
0x103: frame_gpio_obj_group_bin_0163 (RW)
0x104: frame_gpio_obj_group_bin_0274 (RW)
0x105: frame_gpio_obj_group_bin_0030 (RW)
0x106: frame_gpio_obj_group_bin_0135 (RW)
0x107: frame_gpio_obj_group_bin_0256 (RW)
0x108: frame_gpio_obj_group_bin_0012 (RW)
0x109: frame_gpio_obj_group_bin_0123 (RW)
0x10: frame_gpio_obj_group_bin_0000 (RX)
0x10a: frame_gpio_obj_group_bin_0234 (RW)
0x10b: frame_gpio_obj_group_bin_0345 (RW)
0x10c: frame_gpio_obj_group_bin_0101 (RW)
0x10d: frame_gpio_obj_group_bin_0214 (RW)
0x10e: frame_gpio_obj_group_bin_0324 (RW)
0x10f: frame_gpio_obj_group_bin_0083 (RW)
0x110: frame_gpio_obj_group_bin_0193 (RW)
0x111: frame_gpio_obj_group_bin_0303 (RW)
0x112: frame_gpio_obj_group_bin_0062 (RW)
0x113: frame_gpio_obj_group_bin_0173 (RW)
0x114: frame_gpio_obj_group_bin_0282 (RW)
0x115: frame_gpio_obj_group_bin_0040 (RW)
0x116: frame_gpio_obj_group_bin_0153 (RW)
0x117: frame_gpio_obj_group_bin_0156 (RW)
0x118: frame_gpio_obj_group_bin_0021 (RW)
0x119: frame_gpio_obj_group_bin_0134 (RW)
0x11: frame_gpio_obj_group_bin_0001 (RX)
0x11a: frame_gpio_obj_group_bin_0247 (RW)
0x11b: frame_gpio_obj_group_bin_0003 (RW)
0x11c: frame_gpio_obj_group_bin_0114 (RW)
0x11d: frame_gpio_obj_group_bin_0227 (RW)
0x11e: frame_gpio_obj_group_bin_0337 (RW)
0x11f: frame_gpio_obj_group_bin_0094 (RW)
0x120: frame_gpio_obj_group_bin_0206 (RW)
0x121: frame_gpio_obj_group_bin_0316 (RW)
0x122: frame_gpio_obj_group_bin_0075 (RW)
0x123: frame_gpio_obj_group_bin_0185 (RW)
0x124: frame_gpio_obj_group_bin_0295 (RW)
0x125: frame_gpio_obj_group_bin_0054 (RW)
0x126: frame_gpio_obj_group_bin_0165 (RW)
0x127: frame_gpio_obj_group_bin_0275 (RW)
0x128: frame_gpio_obj_group_bin_0032 (RW)
0x129: frame_gpio_obj_group_bin_0145 (RW)
0x12: frame_gpio_obj_group_bin_0240 (RX)
0x12a: frame_gpio_obj_group_bin_0258 (RW)
0x12b: frame_gpio_obj_group_bin_0014 (RW)
0x12c: frame_gpio_obj_group_bin_0125 (RW)
0x12d: frame_gpio_obj_group_bin_0236 (RW)
0x12e: frame_gpio_obj_group_bin_0347 (RW)
0x12f: frame_gpio_obj_group_bin_0103 (RW)
0x130: frame_gpio_obj_group_bin_0216 (RW)
0x131: frame_gpio_obj_group_bin_0326 (RW)
0x132: frame_gpio_obj_group_bin_0085 (RW)
0x133: frame_gpio_obj_group_bin_0195 (RW)
0x134: frame_gpio_obj_group_bin_0305 (RW)
0x135: frame_gpio_obj_group_bin_0064 (RW)
0x136: frame_gpio_obj_group_bin_0175 (RW)
0x138: frame_gpio_obj_group_bin_0042 (RW)
0x13: frame_gpio_obj_group_bin_0351 (RX)
0x13b: frame_gpio_obj_group_bin_0024 (RW)
0x13e: frame_gpio_obj_group_bin_0004 (RW)
0x141: frame_gpio_obj_group_bin_0339 (RW)
0x144: frame_gpio_obj_group_bin_0318 (RW)
0x147: frame_gpio_obj_group_bin_0297 (RW)
0x14: frame_gpio_obj_group_bin_0107 (RX)
0x14a: frame_gpio_obj_group_bin_0277 (RW)
0x14d: frame_gpio_obj_group_bin_0260 (RW)
0x150: frame_gpio_obj_group_bin_0238 (RW)
0x151: frame_gpio_obj_group_bin_0349 (RW)
0x152: frame_gpio_obj_group_bin_0105 (RW)
0x153: frame_gpio_obj_group_bin_0218 (RW)
0x156: frame_gpio_obj_group_bin_0197 (RW)
0x157: frame_gpio_obj_group_bin_0307 (RW)
0x158: frame_gpio_obj_group_bin_0066 (RW)
0x159: frame_gpio_obj_group_bin_0177 (RW)
0x15: frame_gpio_obj_group_bin_0220 (RX)
0x15c: frame_gpio_obj_group_bin_0158 (RW)
0x15d: frame_gpio_obj_group_bin_0270 (RW)
0x15e: frame_gpio_obj_group_bin_0310 (RW)
0x15f: frame_gpio_obj_group_bin_0139 (RW)
0x162: frame_gpio_obj_group_bin_0118 (RW)
0x163: frame_gpio_obj_group_bin_0068 (RW)
0x164: frame_gpio_obj_group_bin_0341 (RW)
0x165: frame_gpio_obj_group_bin_0097 (RW)
0x168: frame_gpio_obj_group_bin_0079 (RW)
0x169: frame_gpio_obj_group_bin_0189 (RW)
0x16: frame_gpio_obj_group_bin_0330 (RX)
0x16a: frame_gpio_obj_group_bin_0299 (RW)
0x16b: frame_gpio_obj_group_bin_0058 (RW)
0x16e: frame_gpio_obj_group_bin_0036 (RW)
0x16f: frame_gpio_obj_group_bin_0149 (RW)
0x170: frame_gpio_obj_group_bin_0262 (RW)
0x171: frame_gpio_obj_group_bin_0018 (RW)
0x174: frame_gpio_obj_group_bin_0352 (RW)
0x175: frame_gpio_obj_group_bin_0108 (RW)
0x176: frame_gpio_obj_group_bin_0221 (RW)
0x177: frame_gpio_obj_group_bin_0331 (RW)
0x17: frame_gpio_obj_group_bin_0089 (RX)
0x17a: frame_gpio_obj_group_bin_0311 (RW)
0x17b: frame_gpio_obj_group_bin_0070 (RW)
0x17c: frame_gpio_obj_group_bin_0180 (RW)
0x17d: frame_gpio_obj_group_bin_0290 (RW)
0x18: frame_gpio_obj_group_bin_0199 (RX)
0x19: frame_gpio_obj_group_bin_0309 (RX)
0x1a: frame_gpio_obj_group_bin_0069 (RX)
0x1b: frame_gpio_obj_group_bin_0246 (RX)
0x1c: frame_gpio_obj_group_bin_0289 (RX)
0x1d: frame_gpio_obj_group_bin_0047 (RX)
0x1e: frame_gpio_obj_group_bin_0160 (RX)
0x1f: frame_gpio_obj_group_bin_0334 (RX)
0x20: frame_gpio_obj_group_bin_0027 (RX)
0x21: frame_gpio_obj_group_bin_0141 (RX)
0x22: frame_gpio_obj_group_bin_0253 (RX)
0x23: frame_gpio_obj_group_bin_0009 (RX)
0x24: frame_gpio_obj_group_bin_0120 (RX)
0x34: frame_gpio_obj_group_bin_0131 (RW)
0x35: frame_gpio_obj_group_bin_0243 (RW)
0x36: frame_gpio_obj_group_bin_0354 (RW)
0x37: frame_gpio_obj_group_bin_0110 (RW)
0x38: frame_gpio_obj_group_bin_0178 (RW)
0x39: frame_gpio_obj_group_bin_0333 (RW)
0x3a: frame_gpio_obj_group_bin_0224 (RW)
0x3b: frame_gpio_obj_group_bin_0203 (RW)
0x3c: frame_gpio_obj_group_bin_0313 (RW)
0x3d: frame_gpio_obj_group_bin_0072 (RW)
0x3e: frame_gpio_obj_group_bin_0182 (RW)
0x3f: frame_gpio_obj_group_bin_0292 (RW)
0x40: frame_gpio_obj_group_bin_0051 (RW)
0x41: frame_gpio_obj_group_bin_0162 (RW)
0x42: frame_gpio_obj_group_bin_0273 (RW)
0x43: frame_gpio_obj_group_bin_0029 (RW)
0x44: frame_gpio_obj_group_bin_0143 (RW)
0x45: frame_gpio_obj_group_bin_0255 (RW)
0x46: frame_gpio_obj_group_bin_0011 (RW)
0x47: frame_gpio_obj_group_bin_0122 (RW)
0x48: frame_gpio_obj_group_bin_0233 (RW)
0x49: frame_gpio_obj_group_bin_0344 (RW)
0x4a: frame_gpio_obj_group_bin_0100 (RW)
0x4b: frame_gpio_obj_group_bin_0213 (RW)
0x4c: frame_gpio_obj_group_bin_0323 (RW)
0x4d: frame_gpio_obj_group_bin_0082 (RW)
0x4e: frame_gpio_obj_group_bin_0192 (RW)
0x4f: frame_gpio_obj_group_bin_0302 (RW)
0x50: frame_gpio_obj_group_bin_0061 (RW)
0x51: frame_gpio_obj_group_bin_0172 (RW)
0x52: frame_gpio_obj_group_bin_0281 (RW)
0x53: frame_gpio_obj_group_bin_0039 (RW)
0x54: frame_gpio_obj_group_bin_0152 (RW)
0x55: frame_gpio_obj_group_bin_0265 (RW)
0x56: frame_gpio_obj_group_bin_0020 (RW)
0x57: frame_gpio_obj_group_bin_0133 (RW)
0x58: frame_gpio_obj_group_bin_0245 (RW)
0x59: frame_gpio_obj_group_bin_0201 (RW)
0x5a: frame_gpio_obj_group_bin_0113 (RW)
0x5b: frame_gpio_obj_group_bin_0226 (RW)
0x5c: frame_gpio_obj_group_bin_0336 (RW)
0x5d: frame_gpio_obj_group_bin_0286 (RW)
0x5e: frame_gpio_obj_group_bin_0205 (RW)
0x5f: frame_gpio_obj_group_bin_0315 (RW)
0x60: frame_gpio_obj_group_bin_0074 (RW)
0x61: frame_gpio_obj_group_bin_0184 (RW)
0x62: frame_gpio_obj_group_bin_0294 (RW)
0x63: frame_gpio_obj_group_bin_0053 (RW)
0x64: frame_gpio_obj_group_bin_0164 (RW)
0x65: frame_gpio_obj_group_bin_0112 (RW)
0x66: frame_gpio_obj_group_bin_0031 (RW)
0x67: frame_gpio_obj_group_bin_0144 (RW)
0x68: frame_gpio_obj_group_bin_0257 (RW)
0x69: frame_gpio_obj_group_bin_0013 (RW)
0x6a: frame_gpio_obj_group_bin_0124 (RW)
0x6b: frame_gpio_obj_group_bin_0235 (RW)
0x6c: frame_gpio_obj_group_bin_0346 (RW)
0x6d: frame_gpio_obj_group_bin_0102 (RW)
0x6e: frame_gpio_obj_group_bin_0215 (RW)
0x6f: frame_gpio_obj_group_bin_0325 (RW)
0x70: frame_gpio_obj_group_bin_0084 (RW)
0x71: frame_gpio_obj_group_bin_0194 (RW)
0x72: frame_gpio_obj_group_bin_0304 (RW)
0x73: frame_gpio_obj_group_bin_0063 (RW)
0x74: frame_gpio_obj_group_bin_0174 (RW)
0x75: frame_gpio_obj_group_bin_0283 (RW)
0x76: frame_gpio_obj_group_bin_0041 (RW)
0x77: frame_gpio_obj_group_bin_0154 (RW)
0x78: frame_gpio_obj_group_bin_0266 (RW)
0x79: frame_gpio_obj_group_bin_0022 (RW)
0x7a: frame_gpio_obj_group_bin_0136 (RW)
0x7b: frame_gpio_obj_group_bin_0248 (RW)
0x7c: frame_gpio_obj_group_bin_0267 (RW)
0x7d: frame_gpio_obj_group_bin_0115 (RW)
0x7e: frame_gpio_obj_group_bin_0228 (RW)
0x7f: frame_gpio_obj_group_bin_0338 (RW)
0x80: frame_gpio_obj_group_bin_0002 (RW)
0x81: frame_gpio_obj_group_bin_0207 (RW)
0x82: frame_gpio_obj_group_bin_0317 (RW)
0x83: frame_gpio_obj_group_bin_0076 (RW)
0x84: frame_gpio_obj_group_bin_0186 (RW)
0x85: frame_gpio_obj_group_bin_0296 (RW)
0x86: frame_gpio_obj_group_bin_0055 (RW)
0x87: frame_gpio_obj_group_bin_0166 (RW)
0x88: frame_gpio_obj_group_bin_0276 (RW)
0x89: frame_gpio_obj_group_bin_0033 (RW)
0x8a: frame_gpio_obj_group_bin_0146 (RW)
0x8b: frame_gpio_obj_group_bin_0259 (RW)
0x8c: frame_gpio_obj_group_bin_0015 (RW)
0x8d: frame_gpio_obj_group_bin_0126 (RW)
0x8e: frame_gpio_obj_group_bin_0237 (RW)
0x8f: frame_gpio_obj_group_bin_0348 (RW)
0x90: frame_gpio_obj_group_bin_0104 (RW)
0x91: frame_gpio_obj_group_bin_0217 (RW)
0x92: frame_gpio_obj_group_bin_0327 (RW)
0x93: frame_gpio_obj_group_bin_0086 (RW)
0x94: frame_gpio_obj_group_bin_0196 (RW)
0x95: frame_gpio_obj_group_bin_0306 (RW)
0x96: frame_gpio_obj_group_bin_0065 (RW)
0x97: frame_gpio_obj_group_bin_0176 (RW)
0x98: frame_gpio_obj_group_bin_0285 (RW)
0x99: frame_gpio_obj_group_bin_0043 (RW)
0x9a: frame_gpio_obj_group_bin_0157 (RW)
0x9b: frame_gpio_obj_group_bin_0269 (RW)
0x9c: frame_gpio_obj_group_bin_0025 (RW)
0x9d: frame_gpio_obj_group_bin_0138 (RW)
0x9e: frame_gpio_obj_group_bin_0250 (RW)
0x9f: frame_gpio_obj_group_bin_0005 (RW)
0xa0: frame_gpio_obj_group_bin_0117 (RW)
0xa1: frame_gpio_obj_group_bin_0230 (RW)
0xa2: frame_gpio_obj_group_bin_0340 (RW)
0xa3: frame_gpio_obj_group_bin_0096 (RW)
0xa4: frame_gpio_obj_group_bin_0209 (RW)
0xa5: frame_gpio_obj_group_bin_0319 (RW)
0xa6: frame_gpio_obj_group_bin_0078 (RW)
0xa7: frame_gpio_obj_group_bin_0188 (RW)
0xa8: frame_gpio_obj_group_bin_0298 (RW)
0xa9: frame_gpio_obj_group_bin_0057 (RW)
0xaa: frame_gpio_obj_group_bin_0168 (RW)
0xab: frame_gpio_obj_group_bin_0278 (RW)
0xac: frame_gpio_obj_group_bin_0035 (RW)
0xad: frame_gpio_obj_group_bin_0148 (RW)
0xae: frame_gpio_obj_group_bin_0261 (RW)
0xaf: frame_gpio_obj_group_bin_0017 (RW)
0xb0: frame_gpio_obj_group_bin_0128 (RW)
0xb1: frame_gpio_obj_group_bin_0239 (RW)
0xb2: frame_gpio_obj_group_bin_0350 (RW)
0xb3: frame_gpio_obj_group_bin_0106 (RW)
0xb4: frame_gpio_obj_group_bin_0219 (RW)
0xb5: frame_gpio_obj_group_bin_0329 (RW)
0xb6: frame_gpio_obj_group_bin_0088 (RW)
0xb7: frame_gpio_obj_group_bin_0198 (RW)
0xb8: frame_gpio_obj_group_bin_0308 (RW)
0xb9: frame_gpio_obj_group_bin_0067 (RW)
0xba: frame_gpio_obj_group_bin_0179 (RW)
0xbb: frame_gpio_obj_group_bin_0288 (RW)
0xbc: frame_gpio_obj_group_bin_0046 (RW)
0xbd: frame_gpio_obj_group_bin_0159 (RW)
0xbe: frame_gpio_obj_group_bin_0271 (RW)
0xbf: frame_gpio_obj_group_bin_0026 (RW)
0xc0: frame_gpio_obj_group_bin_0140 (RW)
0xc1: frame_gpio_obj_group_bin_0252 (RW)
0xc2: frame_gpio_obj_group_bin_0008 (RW)
0xc3: frame_gpio_obj_group_bin_0119 (RW)
0xc4: frame_gpio_obj_group_bin_0092 (RW)
0xc5: frame_gpio_obj_group_bin_0342 (RW)
0xc6: frame_gpio_obj_group_bin_0098 (RW)
0xc7: frame_gpio_obj_group_bin_0211 (RW)
0xc8: frame_gpio_obj_group_bin_0321 (RW)
0xc9: frame_gpio_obj_group_bin_0080 (RW)
0xca: frame_gpio_obj_group_bin_0190 (RW)
0xcb: frame_gpio_obj_group_bin_0300 (RW)
0xcc: frame_gpio_obj_group_bin_0059 (RW)
0xcd: frame_gpio_obj_group_bin_0170 (RW)
0xce: frame_gpio_obj_group_bin_0280 (RW)
0xcf: frame_gpio_obj_group_bin_0037 (RW)
0xd0: frame_gpio_obj_group_bin_0150 (RW)
0xd1: frame_gpio_obj_group_bin_0263 (RW)
0xd2: frame_gpio_obj_group_bin_0044 (RW)
0xd3: frame_gpio_obj_group_bin_0130 (RW)
0xd4: frame_gpio_obj_group_bin_0242 (RW)
0xd5: frame_gpio_obj_group_bin_0353 (RW)
0xd6: frame_gpio_obj_group_bin_0109 (RW)
0xd7: frame_gpio_obj_group_bin_0222 (RW)
0xd8: frame_gpio_obj_group_bin_0332 (RW)
0xd9: frame_gpio_obj_group_bin_0091 (RW)
0xda: frame_gpio_obj_group_bin_0202 (RW)
0xdb: frame_gpio_obj_group_bin_0312 (RW)
0xdc: frame_gpio_obj_group_bin_0071 (RW)
0xdd: frame_gpio_obj_group_bin_0181 (RW)
0xde: frame_gpio_obj_group_bin_0291 (RW)
0xdf: frame_gpio_obj_group_bin_0049 (RW)
0xe0: frame_gpio_obj_group_bin_0161 (RW)
0xe1: frame_gpio_obj_group_bin_0272 (RW)
0xe2: frame_gpio_obj_group_bin_0028 (RW)
0xe3: frame_gpio_obj_group_bin_0142 (RW)
0xe4: frame_gpio_obj_group_bin_0254 (RW)
0xe5: frame_gpio_obj_group_bin_0010 (RW)
0xe6: frame_gpio_obj_group_bin_0121 (RW)
0xe7: frame_gpio_obj_group_bin_0231 (RW)
0xe8: frame_gpio_obj_group_bin_0343 (RW)
0xe9: frame_gpio_obj_group_bin_0099 (RW)
0xea: frame_gpio_obj_group_bin_0212 (RW)
0xeb: frame_gpio_obj_group_bin_0322 (RW)
0xec: frame_gpio_obj_group_bin_0081 (RW)
0xed: frame_gpio_obj_group_bin_0191 (RW)
0xee: frame_gpio_obj_group_bin_0301 (RW)
0xef: frame_gpio_obj_group_bin_0060 (RW)
0xf0: frame_gpio_obj_group_bin_0171 (RW)
0xf1: frame_gpio_obj_group_bin_0023 (RW)
0xf2: frame_gpio_obj_group_bin_0038 (RW)
0xf3: frame_gpio_obj_group_bin_0151 (RW)
0xf4: frame_gpio_obj_group_bin_0264 (RW)
0xf5: frame_gpio_obj_group_bin_0019 (RW)
0xf6: frame_gpio_obj_group_bin_0132 (RW)
0xf7: frame_gpio_obj_group_bin_0244 (RW)
0xf8: frame_gpio_obj_group_bin_0355 (RW)
0xf9: frame_gpio_obj_group_bin_0111 (RW)
0xfa: frame_gpio_obj_group_bin_0225 (RW)
0xfb: frame_gpio_obj_group_bin_0335 (RW)
0xfc: frame_gpio_obj_group_bin_0093 (RW)
0xfd: frame_gpio_obj_group_bin_0204 (RW)
0xfe: frame_gpio_obj_group_bin_0314 (RW)
0xff: frame_gpio_obj_group_bin_0073 (RW)
}
pt_gpio_obj_group_bin_0007 {
0x0: frame_gpio_obj_group_bin_0006 (RW, uncached)
0x100: frame_gpio_obj_group_bin_0223 (RW, uncached)
}
pt_gpio_obj_group_bin_0052 {
0x0: frame_gpio_obj_group_bin_0050 (RW, uncached)
0x100: frame_gpio_obj_group_bin_0232 (RW, uncached)
}
pt_pilot_obj_group_bin_0000 {
0x100: frame_pilot_obj_group_bin_0116 (RW)
0x101: frame_pilot_obj_group_bin_0211 (RW)
0x102: frame_pilot_obj_group_bin_0301 (RW)
0x103: frame_pilot_obj_group_bin_0074 (RW)
0x104: frame_pilot_obj_group_bin_0167 (RW)
0x105: frame_pilot_obj_group_bin_0259 (RW)
0x106: frame_pilot_obj_group_bin_0033 (RW)
0x107: frame_pilot_obj_group_bin_0123 (RW)
0x108: frame_pilot_obj_group_bin_0217 (RW)
0x109: frame_pilot_obj_group_bin_0308 (RW)
0x10: frame_pilot_obj_group_bin_0000 (RX)
0x10a: frame_pilot_obj_group_bin_0081 (RW)
0x10b: frame_pilot_obj_group_bin_0175 (RW)
0x10c: frame_pilot_obj_group_bin_0265 (RW)
0x10d: frame_pilot_obj_group_bin_0039 (RW)
0x10e: frame_pilot_obj_group_bin_0130 (RW)
0x10f: frame_pilot_obj_group_bin_0224 (RW)
0x110: frame_pilot_obj_group_bin_0314 (RW)
0x111: frame_pilot_obj_group_bin_0089 (RW)
0x112: frame_pilot_obj_group_bin_0182 (RW)
0x113: frame_pilot_obj_group_bin_0273 (RW)
0x114: frame_pilot_obj_group_bin_0045 (RW)
0x115: frame_pilot_obj_group_bin_0138 (RW)
0x116: frame_pilot_obj_group_bin_0232 (RW)
0x117: frame_pilot_obj_group_bin_0006 (RW)
0x118: frame_pilot_obj_group_bin_0178 (RW)
0x119: frame_pilot_obj_group_bin_0168 (RW)
0x11: frame_pilot_obj_group_bin_0001 (RX)
0x11a: frame_pilot_obj_group_bin_0075 (RW)
0x11b: frame_pilot_obj_group_bin_0283 (RW)
0x11c: frame_pilot_obj_group_bin_0106 (RW)
0x11d: frame_pilot_obj_group_bin_0251 (RW)
0x11e: frame_pilot_obj_group_bin_0072 (RW)
0x11f: frame_pilot_obj_group_bin_0215 (RW)
0x120: frame_pilot_obj_group_bin_0201 (RW)
0x121: frame_pilot_obj_group_bin_0060 (RW)
0x122: frame_pilot_obj_group_bin_0158 (RW)
0x123: frame_pilot_obj_group_bin_0147 (RW)
0x124: frame_pilot_obj_group_bin_0250 (RW)
0x125: frame_pilot_obj_group_bin_0112 (RW)
0x126: frame_pilot_obj_group_bin_0254 (RW)
0x127: frame_pilot_obj_group_bin_0077 (RW)
0x128: frame_pilot_obj_group_bin_0299 (RW)
0x129: frame_pilot_obj_group_bin_0234 (RW)
0x12: frame_pilot_obj_group_bin_0223 (RX)
0x12a: frame_pilot_obj_group_bin_0165 (RW)
0x12b: frame_pilot_obj_group_bin_0257 (RW)
0x12c: frame_pilot_obj_group_bin_0031 (RW)
0x12d: frame_pilot_obj_group_bin_0121 (RW)
0x12e: frame_pilot_obj_group_bin_0220 (RW)
0x12f: frame_pilot_obj_group_bin_0306 (RW)
0x130: frame_pilot_obj_group_bin_0079 (RW)
0x131: frame_pilot_obj_group_bin_0191 (RW)
0x132: frame_pilot_obj_group_bin_0050 (RW)
0x133: frame_pilot_obj_group_bin_0196 (RW)
0x134: frame_pilot_obj_group_bin_0086 (RW)
0x135: frame_pilot_obj_group_bin_0159 (RW)
0x136: frame_pilot_obj_group_bin_0231 (RW)
0x137: frame_pilot_obj_group_bin_0087 (RW)
0x138: frame_pilot_obj_group_bin_0268 (RW)
0x139: frame_pilot_obj_group_bin_0144 (RW)
0x13: frame_pilot_obj_group_bin_0305 (RX)
0x13a: frame_pilot_obj_group_bin_0235 (RW)
0x13b: frame_pilot_obj_group_bin_0056 (RW)
0x13c: frame_pilot_obj_group_bin_0202 (RW)
0x13d: frame_pilot_obj_group_bin_0025 (RW)
0x13f: frame_pilot_obj_group_bin_0260 (RW)
0x142: frame_pilot_obj_group_bin_0096 (RW)
0x145: frame_pilot_obj_group_bin_0207 (RW)
0x148: frame_pilot_obj_group_bin_0303 (RW)
0x149: frame_pilot_obj_group_bin_0154 (RW)
0x14: frame_pilot_obj_group_bin_0068 (RX)
0x14a: frame_pilot_obj_group_bin_0127 (RW)
0x14b: frame_pilot_obj_group_bin_0022 (RW)
0x14e: frame_pilot_obj_group_bin_0296 (RW)
0x14f: frame_pilot_obj_group_bin_0172 (RW)
0x150: frame_pilot_obj_group_bin_0180 (RW)
0x151: frame_pilot_obj_group_bin_0015 (RW)
0x154: frame_pilot_obj_group_bin_0108 (RW)
0x155: frame_pilot_obj_group_bin_0304 (RW)
0x156: frame_pilot_obj_group_bin_0054 (RW)
0x157: frame_pilot_obj_group_bin_0170 (RW)
0x159: frame_uart_gcs_group_bin_0170 (RWX)
0x15: frame_pilot_obj_group_bin_0151 (RX)
0x15a: frame_pilot_obj_group_bin_0009 (RWX)
0x16: frame_pilot_obj_group_bin_0233 (RX)
0x17: frame_pilot_obj_group_bin_0313 (RX)
0x18: frame_pilot_obj_group_bin_0078 (RX)
0x19: frame_pilot_obj_group_bin_0161 (RX)
0x1a: frame_pilot_obj_group_bin_0162 (RX)
0x1b: frame_pilot_obj_group_bin_0007 (RX)
0x1c: frame_pilot_obj_group_bin_0004 (RX)
0x1d: frame_pilot_obj_group_bin_0171 (RX)
0x1e: frame_pilot_obj_group_bin_0253 (RX)
0x1f: frame_pilot_obj_group_bin_0018 (RX)
0x20: frame_pilot_obj_group_bin_0097 (RX)
0x21: frame_pilot_obj_group_bin_0181 (RX)
0x22: frame_pilot_obj_group_bin_0262 (RX)
0x23: frame_pilot_obj_group_bin_0027 (RX)
0x24: frame_pilot_obj_group_bin_0107 (RX)
0x25: frame_pilot_obj_group_bin_0192 (RX)
0x26: frame_pilot_obj_group_bin_0272 (RX)
0x27: frame_pilot_obj_group_bin_0036 (RX)
0x28: frame_pilot_obj_group_bin_0117 (RX)
0x29: frame_pilot_obj_group_bin_0203 (RX)
0x39: frame_pilot_obj_group_bin_0082 (RW)
0x3a: frame_pilot_obj_group_bin_0005 (RW)
0x3b: frame_pilot_obj_group_bin_0085 (RW)
0x3c: frame_pilot_obj_group_bin_0169 (RW)
0x3d: frame_pilot_obj_group_bin_0252 (RW)
0x3e: frame_pilot_obj_group_bin_0016 (RW)
0x3f: frame_pilot_obj_group_bin_0094 (RW)
0x40: frame_pilot_obj_group_bin_0179 (RW)
0x41: frame_pilot_obj_group_bin_0261 (RW)
0x42: frame_pilot_obj_group_bin_0026 (RW)
0x43: frame_pilot_obj_group_bin_0105 (RW)
0x44: frame_pilot_obj_group_bin_0189 (RW)
0x45: frame_pilot_obj_group_bin_0269 (RW)
0x46: frame_pilot_obj_group_bin_0034 (RW)
0x47: frame_pilot_obj_group_bin_0115 (RW)
0x48: frame_pilot_obj_group_bin_0200 (RW)
0x49: frame_pilot_obj_group_bin_0279 (RW)
0x4a: frame_pilot_obj_group_bin_0042 (RW)
0x4b: frame_pilot_obj_group_bin_0124 (RW)
0x4c: frame_pilot_obj_group_bin_0210 (RW)
0x4d: frame_pilot_obj_group_bin_0291 (RW)
0x4e: frame_pilot_obj_group_bin_0052 (RW)
0x4f: frame_pilot_obj_group_bin_0135 (RW)
0x50: frame_pilot_obj_group_bin_0218 (RW)
0x51: frame_pilot_obj_group_bin_0300 (RW)
0x52: frame_pilot_obj_group_bin_0064 (RW)
0x53: frame_pilot_obj_group_bin_0145 (RW)
0x54: frame_pilot_obj_group_bin_0228 (RW)
0x55: frame_pilot_obj_group_bin_0309 (RW)
0x56: frame_pilot_obj_group_bin_0073 (RW)
0x57: frame_pilot_obj_group_bin_0155 (RW)
0x58: frame_pilot_obj_group_bin_0239 (RW)
0x59: frame_pilot_obj_group_bin_0002 (RW)
0x5a: frame_pilot_obj_group_bin_0083 (RW)
0x5b: frame_pilot_obj_group_bin_0166 (RW)
0x5c: frame_pilot_obj_group_bin_0249 (RW)
0x5d: frame_pilot_obj_group_bin_0013 (RW)
0x5e: frame_pilot_obj_group_bin_0092 (RW)
0x5f: frame_pilot_obj_group_bin_0176 (RW)
0x60: frame_pilot_obj_group_bin_0258 (RW)
0x61: frame_pilot_obj_group_bin_0023 (RW)
0x62: frame_pilot_obj_group_bin_0102 (RW)
0x63: frame_pilot_obj_group_bin_0186 (RW)
0x64: frame_pilot_obj_group_bin_0266 (RW)
0x65: frame_pilot_obj_group_bin_0032 (RW)
0x66: frame_pilot_obj_group_bin_0113 (RW)
0x67: frame_pilot_obj_group_bin_0244 (RW)
0x68: frame_pilot_obj_group_bin_0277 (RW)
0x69: frame_pilot_obj_group_bin_0040 (RW)
0x6a: frame_pilot_obj_group_bin_0122 (RW)
0x6b: frame_pilot_obj_group_bin_0208 (RW)
0x6c: frame_pilot_obj_group_bin_0288 (RW)
0x6d: frame_pilot_obj_group_bin_0049 (RW)
0x6e: frame_pilot_obj_group_bin_0132 (RW)
0x6f: frame_pilot_obj_group_bin_0216 (RW)
0x70: frame_pilot_obj_group_bin_0297 (RW)
0x71: frame_pilot_obj_group_bin_0061 (RW)
0x72: frame_pilot_obj_group_bin_0141 (RW)
0x73: frame_pilot_obj_group_bin_0225 (RW)
0x74: frame_pilot_obj_group_bin_0307 (RW)
0x75: frame_pilot_obj_group_bin_0071 (RW)
0x76: frame_pilot_obj_group_bin_0153 (RW)
0x77: frame_pilot_obj_group_bin_0237 (RW)
0x78: frame_pilot_obj_group_bin_0315 (RW)
0x79: frame_pilot_obj_group_bin_0080 (RW)
0x7a: frame_pilot_obj_group_bin_0163 (RW)
0x7b: frame_pilot_obj_group_bin_0247 (RW)
0x7c: frame_pilot_obj_group_bin_0011 (RW)
0x7d: frame_pilot_obj_group_bin_0090 (RW)
0x7e: frame_pilot_obj_group_bin_0174 (RW)
0x7f: frame_pilot_obj_group_bin_0255 (RW)
0x80: frame_pilot_obj_group_bin_0021 (RW)
0x81: frame_pilot_obj_group_bin_0100 (RW)
0x82: frame_pilot_obj_group_bin_0183 (RW)
0x83: frame_pilot_obj_group_bin_0264 (RW)
0x84: frame_pilot_obj_group_bin_0029 (RW)
0x85: frame_pilot_obj_group_bin_0110 (RW)
0x86: frame_pilot_obj_group_bin_0195 (RW)
0x87: frame_pilot_obj_group_bin_0274 (RW)
0x88: frame_pilot_obj_group_bin_0038 (RW)
0x89: frame_pilot_obj_group_bin_0119 (RW)
0x8a: frame_pilot_obj_group_bin_0205 (RW)
0x8b: frame_pilot_obj_group_bin_0285 (RW)
0x8c: frame_pilot_obj_group_bin_0046 (RW)
0x8d: frame_pilot_obj_group_bin_0129 (RW)
0x8e: frame_pilot_obj_group_bin_0214 (RW)
0x8f: frame_pilot_obj_group_bin_0295 (RW)
0x90: frame_pilot_obj_group_bin_0058 (RW)
0x91: frame_pilot_obj_group_bin_0139 (RW)
0x92: frame_pilot_obj_group_bin_0173 (RW)
0x93: frame_pilot_obj_group_bin_0263 (RW)
0x94: frame_pilot_obj_group_bin_0037 (RW)
0x95: frame_pilot_obj_group_bin_0128 (RW)
0x96: frame_pilot_obj_group_bin_0222 (RW)
0x97: frame_pilot_obj_group_bin_0312 (RW)
0x98: frame_pilot_obj_group_bin_0088 (RW)
0x99: frame_pilot_obj_group_bin_0267 (RW)
0x9a: frame_pilot_obj_group_bin_0245 (RW)
0x9b: frame_pilot_obj_group_bin_0044 (RW)
0x9c: frame_pilot_obj_group_bin_0137 (RW)
0x9d: frame_pilot_obj_group_bin_0230 (RW)
0x9e: frame_pilot_obj_group_bin_0024 (RW)
0x9f: frame_pilot_obj_group_bin_0164 (RW)
0xa0: frame_pilot_obj_group_bin_0190 (RW)
0xa1: frame_pilot_obj_group_bin_0280 (RW)
0xa2: frame_pilot_obj_group_bin_0053 (RW)
0xa3: frame_pilot_obj_group_bin_0146 (RW)
0xa4: frame_pilot_obj_group_bin_0240 (RW)
0xa5: frame_pilot_obj_group_bin_0014 (RW)
0xa6: frame_pilot_obj_group_bin_0103 (RW)
0xa7: frame_pilot_obj_group_bin_0199 (RW)
0xa8: frame_pilot_obj_group_bin_0290 (RW)
0xa9: frame_pilot_obj_group_bin_0062 (RW)
0xaa: frame_pilot_obj_group_bin_0282 (RW)
0xab: frame_pilot_obj_group_bin_0248 (RW)
0xac: frame_pilot_obj_group_bin_0126 (RW)
0xad: frame_pilot_obj_group_bin_0212 (RW)
0xae: frame_pilot_obj_group_bin_0293 (RW)
0xaf: frame_pilot_obj_group_bin_0055 (RW)
0xb0: frame_pilot_obj_group_bin_0070 (RW)
0xb1: frame_pilot_obj_group_bin_0221 (RW)
0xb2: frame_pilot_obj_group_bin_0302 (RW)
0xb3: frame_pilot_obj_group_bin_0066 (RW)
0xb4: frame_pilot_obj_group_bin_0148 (RW)
0xb5: frame_pilot_obj_group_bin_0213 (RW)
0xb6: frame_pilot_obj_group_bin_0311 (RW)
0xb7: frame_pilot_obj_group_bin_0076 (RW)
0xb8: frame_pilot_obj_group_bin_0157 (RW)
0xb9: frame_pilot_obj_group_bin_0242 (RW)
0xba: frame_pilot_obj_group_bin_0184 (RW)
0xbb: frame_pilot_obj_group_bin_0008 (RW)
0xbc: frame_pilot_obj_group_bin_0149 (RW)
0xbd: frame_pilot_obj_group_bin_0292 (RW)
0xbe: frame_pilot_obj_group_bin_0114 (RW)
0xbf: frame_pilot_obj_group_bin_0256 (RW)
0xc0: frame_pilot_obj_group_bin_0270 (RW)
0xc1: frame_pilot_obj_group_bin_0043 (RW)
0xc2: frame_pilot_obj_group_bin_0136 (RW)
0xc3: frame_pilot_obj_group_bin_0229 (RW)
0xc4: frame_pilot_obj_group_bin_0003 (RW)
0xc5: frame_pilot_obj_group_bin_0093 (RW)
0xc6: frame_pilot_obj_group_bin_0187 (RW)
0xc7: frame_pilot_obj_group_bin_0278 (RW)
0xc8: frame_pilot_obj_group_bin_0051 (RW)
0xc9: frame_pilot_obj_group_bin_0143 (RW)
0xca: frame_pilot_obj_group_bin_0238 (RW)
0xcb: frame_pilot_obj_group_bin_0012 (RW)
0xcc: frame_pilot_obj_group_bin_0101 (RW)
0xcd: frame_pilot_obj_group_bin_0197 (RW)
0xce: frame_pilot_obj_group_bin_0286 (RW)
0xcf: frame_pilot_obj_group_bin_0059 (RW)
0xd0: frame_pilot_obj_group_bin_0152 (RW)
0xd1: frame_pilot_obj_group_bin_0246 (RW)
0xd2: frame_pilot_obj_group_bin_0020 (RW)
0xd3: frame_pilot_obj_group_bin_0109 (RW)
0xd4: frame_pilot_obj_group_bin_0204 (RW)
0xd5: frame_pilot_obj_group_bin_0294 (RW)
0xd6: frame_pilot_obj_group_bin_0067 (RW)
0xd7: frame_pilot_obj_group_bin_0160 (RW)
0xd8: frame_pilot_obj_group_bin_0310 (RW)
0xd9: frame_pilot_obj_group_bin_0133 (RW)
0xda: frame_pilot_obj_group_bin_0275 (RW)
0xdb: frame_pilot_obj_group_bin_0098 (RW)
0xdc: frame_pilot_obj_group_bin_0243 (RW)
0xdd: frame_pilot_obj_group_bin_0065 (RW)
0xde: frame_pilot_obj_group_bin_0209 (RW)
0xdf: frame_pilot_obj_group_bin_0030 (RW)
0xe0: frame_pilot_obj_group_bin_0035 (RW)
0xe1: frame_pilot_obj_group_bin_0125 (RW)
0xe2: frame_pilot_obj_group_bin_0219 (RW)
0xe3: frame_pilot_obj_group_bin_0281 (RW)
0xe4: frame_pilot_obj_group_bin_0084 (RW)
0xe5: frame_pilot_obj_group_bin_0177 (RW)
0xe6: frame_pilot_obj_group_bin_0069 (RW)
0xe7: frame_pilot_obj_group_bin_0198 (RW)
0xe8: frame_pilot_obj_group_bin_0134 (RW)
0xe9: frame_pilot_obj_group_bin_0227 (RW)
0xea: frame_pilot_obj_group_bin_0095 (RW)
0xeb: frame_pilot_obj_group_bin_0091 (RW)
0xec: frame_pilot_obj_group_bin_0185 (RW)
0xed: frame_pilot_obj_group_bin_0276 (RW)
0xee: frame_pilot_obj_group_bin_0048 (RW)
0xef: frame_pilot_obj_group_bin_0140 (RW)
0xf0: frame_pilot_obj_group_bin_0236 (RW)
0xf1: frame_pilot_obj_group_bin_0010 (RW)
0xf2: frame_pilot_obj_group_bin_0099 (RW)
0xf3: frame_pilot_obj_group_bin_0194 (RW)
0xf4: frame_pilot_obj_group_bin_0284 (RW)
0xf5: frame_pilot_obj_group_bin_0057 (RW)
0xf6: frame_pilot_obj_group_bin_0150 (RW)
0xf7: frame_pilot_obj_group_bin_0019 (RW)
0xf8: frame_pilot_obj_group_bin_0104 (RW)
0xf9: frame_pilot_obj_group_bin_0226 (RW)
0xfa: frame_pilot_obj_group_bin_0047 (RW)
0xfb: frame_pilot_obj_group_bin_0193 (RW)
0xfc: frame_pilot_obj_group_bin_0017 (RW)
0xfd: frame_pilot_obj_group_bin_0156 (RW)
0xfe: frame_pilot_obj_group_bin_0298 (RW)
0xff: frame_pilot_obj_group_bin_0120 (RW)
}
pt_pwm_obj_group_bin_0000 {
0x100: frame_pwm_obj_group_bin_0122 (RW)
0x101: frame_pwm_obj_group_bin_0220 (RW)
0x102: frame_pwm_obj_group_bin_0319 (RW)
0x103: frame_pwm_obj_group_bin_0077 (RW)
0x104: frame_pwm_obj_group_bin_0175 (RW)
0x105: frame_pwm_obj_group_bin_0271 (RW)
0x106: frame_pwm_obj_group_bin_0036 (RW)
0x107: frame_pwm_obj_group_bin_0129 (RW)
0x108: frame_pwm_obj_group_bin_0226 (RW)
0x109: frame_pwm_obj_group_bin_0325 (RW)
0x10: frame_pwm_obj_group_bin_0000 (RX)
0x10a: frame_pwm_obj_group_bin_0085 (RW)
0x10b: frame_pwm_obj_group_bin_0183 (RW)
0x10c: frame_pwm_obj_group_bin_0280 (RW)
0x10d: frame_pwm_obj_group_bin_0042 (RW)
0x10e: frame_pwm_obj_group_bin_0136 (RW)
0x10f: frame_pwm_obj_group_bin_0233 (RW)
0x110: frame_pwm_obj_group_bin_0333 (RW)
0x111: frame_pwm_obj_group_bin_0093 (RW)
0x112: frame_pwm_obj_group_bin_0190 (RW)
0x113: frame_pwm_obj_group_bin_0288 (RW)
0x114: frame_pwm_obj_group_bin_0050 (RW)
0x115: frame_pwm_obj_group_bin_0144 (RW)
0x116: frame_pwm_obj_group_bin_0242 (RW)
0x117: frame_pwm_obj_group_bin_0006 (RW)
0x118: frame_pwm_obj_group_bin_0186 (RW)
0x119: frame_pwm_obj_group_bin_0176 (RW)
0x11: frame_pwm_obj_group_bin_0001 (RX)
0x11a: frame_pwm_obj_group_bin_0078 (RW)
0x11b: frame_pwm_obj_group_bin_0298 (RW)
0x11c: frame_pwm_obj_group_bin_0111 (RW)
0x11d: frame_pwm_obj_group_bin_0262 (RW)
0x11e: frame_pwm_obj_group_bin_0075 (RW)
0x11f: frame_pwm_obj_group_bin_0224 (RW)
0x120: frame_pwm_obj_group_bin_0043 (RW)
0x121: frame_pwm_obj_group_bin_0307 (RW)
0x122: frame_pwm_obj_group_bin_0166 (RW)
0x123: frame_pwm_obj_group_bin_0152 (RW)
0x124: frame_pwm_obj_group_bin_0261 (RW)
0x125: frame_pwm_obj_group_bin_0117 (RW)
0x126: frame_pwm_obj_group_bin_0266 (RW)
0x127: frame_pwm_obj_group_bin_0055 (RW)
0x128: frame_pwm_obj_group_bin_0317 (RW)
0x129: frame_pwm_obj_group_bin_0244 (RW)
0x12: frame_pwm_obj_group_bin_0232 (RX)
0x12a: frame_pwm_obj_group_bin_0173 (RW)
0x12b: frame_pwm_obj_group_bin_0269 (RW)
0x12c: frame_pwm_obj_group_bin_0034 (RW)
0x12d: frame_pwm_obj_group_bin_0127 (RW)
0x12e: frame_pwm_obj_group_bin_0229 (RW)
0x12f: frame_pwm_obj_group_bin_0323 (RW)
0x130: frame_pwm_obj_group_bin_0083 (RW)
0x131: frame_pwm_obj_group_bin_0199 (RW)
0x132: frame_pwm_obj_group_bin_0275 (RW)
0x133: frame_pwm_obj_group_bin_0205 (RW)
0x134: frame_pwm_obj_group_bin_0090 (RW)
0x135: frame_pwm_obj_group_bin_0167 (RW)
0x136: frame_pwm_obj_group_bin_0241 (RW)
0x138: frame_pwm_obj_group_bin_0283 (RW)
0x13: frame_pwm_obj_group_bin_0322 (RX)
0x13b: frame_pwm_obj_group_bin_0061 (RW)
0x13e: frame_pwm_obj_group_bin_0196 (RW)
0x141: frame_pwm_obj_group_bin_0286 (RW)
0x144: frame_pwm_obj_group_bin_0015 (RW)
0x147: frame_pwm_obj_group_bin_0305 (RW)
0x14: frame_pwm_obj_group_bin_0071 (RX)
0x14a: frame_pwm_obj_group_bin_0133 (RW)
0x14b: frame_pwm_obj_group_bin_0024 (RW)
0x14c: frame_pwm_obj_group_bin_0116 (RW)
0x14d: frame_pwm_obj_group_bin_0216 (RW)
0x150: frame_pwm_obj_group_bin_0188 (RW)
0x151: frame_pwm_obj_group_bin_0016 (RW)
0x152: frame_pwm_obj_group_bin_0031 (RW)
0x153: frame_pwm_obj_group_bin_0301 (RW)
0x156: frame_pwm_obj_group_bin_0059 (RW)
0x157: frame_pwm_obj_group_bin_0178 (RW)
0x158: frame_pwm_obj_group_bin_0046 (RW)
0x159: frame_pwm_obj_group_bin_0303 (RW)
0x15: frame_pwm_obj_group_bin_0157 (RX)
0x15c: frame_pwm_obj_group_bin_0308 (RW)
0x15d: frame_pwm_obj_group_bin_0120 (RW)
0x15e: frame_pwm_obj_group_bin_0013 (RW)
0x15f: frame_pwm_obj_group_bin_0082 (RW)
0x162: frame_pwm_obj_group_bin_0200 (RW)
0x163: frame_pwm_obj_group_bin_0017 (RW)
0x164: frame_pwm_obj_group_bin_0162 (RW)
0x165: frame_pwm_obj_group_bin_0314 (RW)
0x168: frame_pwm_obj_group_bin_0326 (RW)
0x169: frame_pwm_obj_group_bin_0312 (RW)
0x16: frame_pwm_obj_group_bin_0243 (RX)
0x16a: frame_pwm_obj_group_bin_0098 (RW)
0x16b: frame_pwm_obj_group_bin_0029 (RW)
0x17: frame_pwm_obj_group_bin_0331 (RX)
0x18: frame_pwm_obj_group_bin_0081 (RX)
0x19: frame_pwm_obj_group_bin_0169 (RX)
0x1a: frame_pwm_obj_group_bin_0170 (RX)
0x1b: frame_pwm_obj_group_bin_0007 (RX)
0x1c: frame_pwm_obj_group_bin_0092 (RX)
0x1d: frame_pwm_obj_group_bin_0179 (RX)
0x1e: frame_pwm_obj_group_bin_0265 (RX)
0x1f: frame_pwm_obj_group_bin_0020 (RX)
0x20: frame_pwm_obj_group_bin_0102 (RX)
0x21: frame_pwm_obj_group_bin_0189 (RX)
0x22: frame_pwm_obj_group_bin_0277 (RX)
0x23: frame_pwm_obj_group_bin_0030 (RX)
0x24: frame_pwm_obj_group_bin_0112 (RX)
0x34: frame_pwm_obj_group_bin_0153 (RW)
0x35: frame_pwm_obj_group_bin_0240 (RW)
0x36: frame_pwm_obj_group_bin_0329 (RW)
0x37: frame_pwm_obj_group_bin_0079 (RW)
0x38: frame_pwm_obj_group_bin_0004 (RW)
0x39: frame_pwm_obj_group_bin_0252 (RW)
0x3a: frame_pwm_obj_group_bin_0005 (RW)
0x3b: frame_pwm_obj_group_bin_0089 (RW)
0x3c: frame_pwm_obj_group_bin_0177 (RW)
0x3d: frame_pwm_obj_group_bin_0086 (RW)
0x3e: frame_pwm_obj_group_bin_0018 (RW)
0x3f: frame_pwm_obj_group_bin_0099 (RW)
0x40: frame_pwm_obj_group_bin_0187 (RW)
0x41: frame_pwm_obj_group_bin_0273 (RW)
0x42: frame_pwm_obj_group_bin_0028 (RW)
0x43: frame_pwm_obj_group_bin_0110 (RW)
0x44: frame_pwm_obj_group_bin_0197 (RW)
0x45: frame_pwm_obj_group_bin_0284 (RW)
0x46: frame_pwm_obj_group_bin_0037 (RW)
0x47: frame_pwm_obj_group_bin_0121 (RW)
0x48: frame_pwm_obj_group_bin_0209 (RW)
0x49: frame_pwm_obj_group_bin_0294 (RW)
0x4a: frame_pwm_obj_group_bin_0047 (RW)
0x4b: frame_pwm_obj_group_bin_0130 (RW)
0x4c: frame_pwm_obj_group_bin_0219 (RW)
0x4d: frame_pwm_obj_group_bin_0306 (RW)
0x4e: frame_pwm_obj_group_bin_0057 (RW)
0x4f: frame_pwm_obj_group_bin_0141 (RW)
0x50: frame_pwm_obj_group_bin_0227 (RW)
0x51: frame_pwm_obj_group_bin_0318 (RW)
0x52: frame_pwm_obj_group_bin_0067 (RW)
0x53: frame_pwm_obj_group_bin_0150 (RW)
0x54: frame_pwm_obj_group_bin_0238 (RW)
0x55: frame_pwm_obj_group_bin_0327 (RW)
0x56: frame_pwm_obj_group_bin_0076 (RW)
0x57: frame_pwm_obj_group_bin_0163 (RW)
0x58: frame_pwm_obj_group_bin_0249 (RW)
0x59: frame_pwm_obj_group_bin_0002 (RW)
0x5a: frame_pwm_obj_group_bin_0087 (RW)
0x5b: frame_pwm_obj_group_bin_0174 (RW)
0x5c: frame_pwm_obj_group_bin_0260 (RW)
0x5d: frame_pwm_obj_group_bin_0014 (RW)
0x5e: frame_pwm_obj_group_bin_0096 (RW)
0x5f: frame_pwm_obj_group_bin_0184 (RW)
0x60: frame_pwm_obj_group_bin_0270 (RW)
0x61: frame_pwm_obj_group_bin_0025 (RW)
0x62: frame_pwm_obj_group_bin_0107 (RW)
0x63: frame_pwm_obj_group_bin_0194 (RW)
0x64: frame_pwm_obj_group_bin_0281 (RW)
0x65: frame_pwm_obj_group_bin_0035 (RW)
0x66: frame_pwm_obj_group_bin_0118 (RW)
0x67: frame_pwm_obj_group_bin_0254 (RW)
0x68: frame_pwm_obj_group_bin_0292 (RW)
0x69: frame_pwm_obj_group_bin_0044 (RW)
0x6a: frame_pwm_obj_group_bin_0128 (RW)
0x6b: frame_pwm_obj_group_bin_0217 (RW)
0x6c: frame_pwm_obj_group_bin_0304 (RW)
0x6d: frame_pwm_obj_group_bin_0054 (RW)
0x6e: frame_pwm_obj_group_bin_0138 (RW)
0x6f: frame_pwm_obj_group_bin_0225 (RW)
0x70: frame_pwm_obj_group_bin_0315 (RW)
0x71: frame_pwm_obj_group_bin_0065 (RW)
0x72: frame_pwm_obj_group_bin_0147 (RW)
0x73: frame_pwm_obj_group_bin_0235 (RW)
0x74: frame_pwm_obj_group_bin_0324 (RW)
0x75: frame_pwm_obj_group_bin_0074 (RW)
0x76: frame_pwm_obj_group_bin_0159 (RW)
0x77: frame_pwm_obj_group_bin_0247 (RW)
0x78: frame_pwm_obj_group_bin_0334 (RW)
0x79: frame_pwm_obj_group_bin_0084 (RW)
0x7a: frame_pwm_obj_group_bin_0171 (RW)
0x7b: frame_pwm_obj_group_bin_0257 (RW)
0x7c: frame_pwm_obj_group_bin_0011 (RW)
0x7d: frame_pwm_obj_group_bin_0094 (RW)
0x7e: frame_pwm_obj_group_bin_0182 (RW)
0x7f: frame_pwm_obj_group_bin_0267 (RW)
0x80: frame_pwm_obj_group_bin_0023 (RW)
0x81: frame_pwm_obj_group_bin_0105 (RW)
0x82: frame_pwm_obj_group_bin_0191 (RW)
0x83: frame_pwm_obj_group_bin_0279 (RW)
0x84: frame_pwm_obj_group_bin_0032 (RW)
0x85: frame_pwm_obj_group_bin_0115 (RW)
0x86: frame_pwm_obj_group_bin_0204 (RW)
0x87: frame_pwm_obj_group_bin_0289 (RW)
0x88: frame_pwm_obj_group_bin_0041 (RW)
0x89: frame_pwm_obj_group_bin_0125 (RW)
0x8a: frame_pwm_obj_group_bin_0215 (RW)
0x8b: frame_pwm_obj_group_bin_0300 (RW)
0x8c: frame_pwm_obj_group_bin_0051 (RW)
0x8d: frame_pwm_obj_group_bin_0135 (RW)
0x8e: frame_pwm_obj_group_bin_0223 (RW)
0x8f: frame_pwm_obj_group_bin_0311 (RW)
0x90: frame_pwm_obj_group_bin_0063 (RW)
0x91: frame_pwm_obj_group_bin_0145 (RW)
0x92: frame_pwm_obj_group_bin_0181 (RW)
0x93: frame_pwm_obj_group_bin_0278 (RW)
0x94: frame_pwm_obj_group_bin_0040 (RW)
0x95: frame_pwm_obj_group_bin_0134 (RW)
0x96: frame_pwm_obj_group_bin_0231 (RW)
0x97: frame_pwm_obj_group_bin_0330 (RW)
0x98: frame_pwm_obj_group_bin_0131 (RW)
0x99: frame_pwm_obj_group_bin_0282 (RW)
0x9a: frame_pwm_obj_group_bin_0255 (RW)
0x9b: frame_pwm_obj_group_bin_0049 (RW)
0x9c: frame_pwm_obj_group_bin_0143 (RW)
0x9d: frame_pwm_obj_group_bin_0210 (RW)
0x9e: frame_pwm_obj_group_bin_0026 (RW)
0x9f: frame_pwm_obj_group_bin_0172 (RW)
0xa0: frame_pwm_obj_group_bin_0198 (RW)
0xa1: frame_pwm_obj_group_bin_0295 (RW)
0xa2: frame_pwm_obj_group_bin_0058 (RW)
0xa3: frame_pwm_obj_group_bin_0151 (RW)
0xa4: frame_pwm_obj_group_bin_0250 (RW)
0xa5: frame_pwm_obj_group_bin_0201 (RW)
0xa6: frame_pwm_obj_group_bin_0287 (RW)
0xa7: frame_pwm_obj_group_bin_0039 (RW)
0xa8: frame_pwm_obj_group_bin_0123 (RW)
0xa9: frame_pwm_obj_group_bin_0213 (RW)
0xaa: frame_pwm_obj_group_bin_0297 (RW)
0xab: frame_pwm_obj_group_bin_0259 (RW)
0xac: frame_pwm_obj_group_bin_0132 (RW)
0xad: frame_pwm_obj_group_bin_0221 (RW)
0xae: frame_pwm_obj_group_bin_0309 (RW)
0xaf: frame_pwm_obj_group_bin_0060 (RW)
0xb0: frame_pwm_obj_group_bin_0073 (RW)
0xb1: frame_pwm_obj_group_bin_0230 (RW)
0xb2: frame_pwm_obj_group_bin_0320 (RW)
0xb3: frame_pwm_obj_group_bin_0069 (RW)
0xb4: frame_pwm_obj_group_bin_0124 (RW)
0xb5: frame_pwm_obj_group_bin_0222 (RW)
0xb6: frame_pwm_obj_group_bin_0321 (RW)
0xb7: frame_pwm_obj_group_bin_0080 (RW)
0xb8: frame_pwm_obj_group_bin_0165 (RW)
0xb9: frame_pwm_obj_group_bin_0045 (RW)
0xba: frame_pwm_obj_group_bin_0192 (RW)
0xbb: frame_pwm_obj_group_bin_0008 (RW)
0xbc: frame_pwm_obj_group_bin_0154 (RW)
0xbd: frame_pwm_obj_group_bin_0263 (RW)
0xbe: frame_pwm_obj_group_bin_0119 (RW)
0xbf: frame_pwm_obj_group_bin_0268 (RW)
0xc0: frame_pwm_obj_group_bin_0285 (RW)
0xc1: frame_pwm_obj_group_bin_0048 (RW)
0xc2: frame_pwm_obj_group_bin_0142 (RW)
0xc3: frame_pwm_obj_group_bin_0239 (RW)
0xc4: frame_pwm_obj_group_bin_0003 (RW)
0xc5: frame_pwm_obj_group_bin_0097 (RW)
0xc6: frame_pwm_obj_group_bin_0195 (RW)
0xc7: frame_pwm_obj_group_bin_0293 (RW)
0xc8: frame_pwm_obj_group_bin_0056 (RW)
0xc9: frame_pwm_obj_group_bin_0148 (RW)
0xca: frame_pwm_obj_group_bin_0248 (RW)
0xcb: frame_pwm_obj_group_bin_0012 (RW)
0xcc: frame_pwm_obj_group_bin_0106 (RW)
0xcd: frame_pwm_obj_group_bin_0206 (RW)
0xce: frame_pwm_obj_group_bin_0302 (RW)
0xcf: frame_pwm_obj_group_bin_0064 (RW)
0xd0: frame_pwm_obj_group_bin_0158 (RW)
0xd1: frame_pwm_obj_group_bin_0256 (RW)
0xd2: frame_pwm_obj_group_bin_0022 (RW)
0xd3: frame_pwm_obj_group_bin_0114 (RW)
0xd4: frame_pwm_obj_group_bin_0214 (RW)
0xd5: frame_pwm_obj_group_bin_0310 (RW)
0xd6: frame_pwm_obj_group_bin_0070 (RW)
0xd7: frame_pwm_obj_group_bin_0168 (RW)
0xd8: frame_pwm_obj_group_bin_0328 (RW)
0xd9: frame_pwm_obj_group_bin_0139 (RW)
0xda: frame_pwm_obj_group_bin_0290 (RW)
0xdb: frame_pwm_obj_group_bin_0103 (RW)
0xdc: frame_pwm_obj_group_bin_0253 (RW)
0xdd: frame_pwm_obj_group_bin_0068 (RW)
0xde: frame_pwm_obj_group_bin_0218 (RW)
0xdf: frame_pwm_obj_group_bin_0033 (RW)
0xe0: frame_pwm_obj_group_bin_0038 (RW)
0xe1: frame_pwm_obj_group_bin_0332 (RW)
0xe2: frame_pwm_obj_group_bin_0228 (RW)
0xe3: frame_pwm_obj_group_bin_0296 (RW)
0xe4: frame_pwm_obj_group_bin_0088 (RW)
0xe5: frame_pwm_obj_group_bin_0185 (RW)
0xe6: frame_pwm_obj_group_bin_0072 (RW)
0xe7: frame_pwm_obj_group_bin_0207 (RW)
0xe8: frame_pwm_obj_group_bin_0140 (RW)
0xe9: frame_pwm_obj_group_bin_0237 (RW)
0xea: frame_pwm_obj_group_bin_0100 (RW)
0xeb: frame_pwm_obj_group_bin_0095 (RW)
0xec: frame_pwm_obj_group_bin_0193 (RW)
0xed: frame_pwm_obj_group_bin_0291 (RW)
0xee: frame_pwm_obj_group_bin_0053 (RW)
0xef: frame_pwm_obj_group_bin_0146 (RW)
0xf0: frame_pwm_obj_group_bin_0246 (RW)
0xf1: frame_pwm_obj_group_bin_0010 (RW)
0xf2: frame_pwm_obj_group_bin_0104 (RW)
0xf3: frame_pwm_obj_group_bin_0203 (RW)
0xf4: frame_pwm_obj_group_bin_0299 (RW)
0xf5: frame_pwm_obj_group_bin_0062 (RW)
0xf6: frame_pwm_obj_group_bin_0156 (RW)
0xf7: frame_pwm_obj_group_bin_0021 (RW)
0xf8: frame_pwm_obj_group_bin_0109 (RW)
0xf9: frame_pwm_obj_group_bin_0236 (RW)
0xfa: frame_pwm_obj_group_bin_0052 (RW)
0xfb: frame_pwm_obj_group_bin_0202 (RW)
0xfc: frame_pwm_obj_group_bin_0019 (RW)
0xfd: frame_pwm_obj_group_bin_0164 (RW)
0xfe: frame_pwm_obj_group_bin_0316 (RW)
0xff: frame_pwm_obj_group_bin_0126 (RW)
}
pt_pwm_obj_group_bin_0259 {
0x0: frame_pwm_obj_group_bin_0258 (RW, uncached)
}
pt_spi_obj_group_bin_0000 {
0x100: frame_spi_obj_group_bin_0116 (RW)
0x101: frame_spi_obj_group_bin_0210 (RW)
0x102: frame_spi_obj_group_bin_0302 (RW)
0x103: frame_spi_obj_group_bin_0074 (RW)
0x104: frame_spi_obj_group_bin_0167 (RW)
0x105: frame_spi_obj_group_bin_0259 (RW)
0x106: frame_spi_obj_group_bin_0033 (RW)
0x107: frame_spi_obj_group_bin_0123 (RW)
0x108: frame_spi_obj_group_bin_0216 (RW)
0x109: frame_spi_obj_group_bin_0308 (RW)
0x10: frame_spi_obj_group_bin_0000 (RX)
0x10a: frame_spi_obj_group_bin_0081 (RW)
0x10b: frame_spi_obj_group_bin_0175 (RW)
0x10c: frame_spi_obj_group_bin_0266 (RW)
0x10d: frame_spi_obj_group_bin_0039 (RW)
0x10e: frame_spi_obj_group_bin_0130 (RW)
0x10f: frame_spi_obj_group_bin_0223 (RW)
0x110: frame_spi_obj_group_bin_0315 (RW)
0x111: frame_spi_obj_group_bin_0089 (RW)
0x112: frame_spi_obj_group_bin_0182 (RW)
0x113: frame_spi_obj_group_bin_0274 (RW)
0x114: frame_spi_obj_group_bin_0047 (RW)
0x115: frame_spi_obj_group_bin_0138 (RW)
0x116: frame_spi_obj_group_bin_0231 (RW)
0x117: frame_spi_obj_group_bin_0006 (RW)
0x118: frame_spi_obj_group_bin_0178 (RW)
0x119: frame_spi_obj_group_bin_0168 (RW)
0x11: frame_spi_obj_group_bin_0001 (RX)
0x11a: frame_spi_obj_group_bin_0075 (RW)
0x11b: frame_spi_obj_group_bin_0284 (RW)
0x11c: frame_spi_obj_group_bin_0106 (RW)
0x11d: frame_spi_obj_group_bin_0250 (RW)
0x11e: frame_spi_obj_group_bin_0072 (RW)
0x11f: frame_spi_obj_group_bin_0214 (RW)
0x120: frame_spi_obj_group_bin_0040 (RW)
0x121: frame_spi_obj_group_bin_0293 (RW)
0x122: frame_spi_obj_group_bin_0158 (RW)
0x123: frame_spi_obj_group_bin_0147 (RW)
0x124: frame_spi_obj_group_bin_0249 (RW)
0x125: frame_spi_obj_group_bin_0112 (RW)
0x126: frame_spi_obj_group_bin_0254 (RW)
0x127: frame_spi_obj_group_bin_0052 (RW)
0x128: frame_spi_obj_group_bin_0300 (RW)
0x129: frame_spi_obj_group_bin_0233 (RW)
0x12: frame_spi_obj_group_bin_0222 (RX)
0x12a: frame_spi_obj_group_bin_0165 (RW)
0x12b: frame_spi_obj_group_bin_0257 (RW)
0x12c: frame_spi_obj_group_bin_0031 (RW)
0x12d: frame_spi_obj_group_bin_0121 (RW)
0x12e: frame_spi_obj_group_bin_0219 (RW)
0x12f: frame_spi_obj_group_bin_0306 (RW)
0x130: frame_spi_obj_group_bin_0079 (RW)
0x131: frame_spi_obj_group_bin_0191 (RW)
0x132: frame_spi_obj_group_bin_0262 (RW)
0x133: frame_spi_obj_group_bin_0196 (RW)
0x134: frame_spi_obj_group_bin_0086 (RW)
0x135: frame_spi_obj_group_bin_0159 (RW)
0x137: frame_spi_obj_group_bin_0087 (RW)
0x13: frame_spi_obj_group_bin_0305 (RX)
0x13a: frame_spi_obj_group_bin_0234 (RW)
0x13d: frame_spi_obj_group_bin_0025 (RW)
0x140: frame_spi_obj_group_bin_0131 (RW)
0x143: frame_spi_obj_group_bin_0239 (RW)
0x144: frame_spi_obj_group_bin_0014 (RW)
0x145: frame_spi_obj_group_bin_0103 (RW)
0x146: frame_spi_obj_group_bin_0199 (RW)
0x149: frame_spi_obj_group_bin_0154 (RW)
0x14: frame_spi_obj_group_bin_0068 (RX)
0x14a: frame_spi_obj_group_bin_0127 (RW)
0x14b: frame_spi_obj_group_bin_0022 (RW)
0x14c: frame_spi_obj_group_bin_0111 (RW)
0x14f: frame_spi_obj_group_bin_0172 (RW)
0x150: frame_spi_obj_group_bin_0180 (RW)
0x151: frame_spi_obj_group_bin_0015 (RW)
0x152: frame_spi_obj_group_bin_0142 (RW)
0x155: frame_spi_obj_group_bin_0252 (RW)
0x156: frame_spi_obj_group_bin_0056 (RW)
0x157: frame_spi_obj_group_bin_0170 (RW)
0x158: frame_spi_obj_group_bin_0043 (RW)
0x15: frame_spi_obj_group_bin_0151 (RX)
0x15a: frame_can_obj_group_bin_0284 (RWX)
0x16: frame_spi_obj_group_bin_0232 (RX)
0x17: frame_spi_obj_group_bin_0313 (RX)
0x18: frame_spi_obj_group_bin_0078 (RX)
0x19: frame_spi_obj_group_bin_0161 (RX)
0x1a: frame_spi_obj_group_bin_0162 (RX)
0x1b: frame_spi_obj_group_bin_0007 (RX)
0x1c: frame_spi_obj_group_bin_0088 (RX)
0x1d: frame_spi_obj_group_bin_0171 (RX)
0x1e: frame_spi_obj_group_bin_0253 (RX)
0x1f: frame_spi_obj_group_bin_0018 (RX)
0x20: frame_spi_obj_group_bin_0097 (RX)
0x21: frame_spi_obj_group_bin_0181 (RX)
0x22: frame_spi_obj_group_bin_0263 (RX)
0x23: frame_spi_obj_group_bin_0027 (RX)
0x33: frame_spi_obj_group_bin_0066 (RW)
0x34: frame_spi_obj_group_bin_0148 (RW)
0x35: frame_spi_obj_group_bin_0229 (RW)
0x36: frame_spi_obj_group_bin_0311 (RW)
0x37: frame_spi_obj_group_bin_0076 (RW)
0x38: frame_spi_obj_group_bin_0004 (RW)
0x39: frame_spi_obj_group_bin_0240 (RW)
0x3a: frame_spi_obj_group_bin_0005 (RW)
0x3b: frame_spi_obj_group_bin_0085 (RW)
0x3c: frame_spi_obj_group_bin_0169 (RW)
0x3d: frame_spi_obj_group_bin_0082 (RW)
0x3e: frame_spi_obj_group_bin_0016 (RW)
0x3f: frame_spi_obj_group_bin_0094 (RW)
0x40: frame_spi_obj_group_bin_0179 (RW)
0x41: frame_spi_obj_group_bin_0261 (RW)
0x42: frame_spi_obj_group_bin_0026 (RW)
0x43: frame_spi_obj_group_bin_0105 (RW)
0x44: frame_spi_obj_group_bin_0189 (RW)
0x45: frame_spi_obj_group_bin_0270 (RW)
0x46: frame_spi_obj_group_bin_0034 (RW)
0x47: frame_spi_obj_group_bin_0115 (RW)
0x48: frame_spi_obj_group_bin_0200 (RW)
0x49: frame_spi_obj_group_bin_0280 (RW)
0x4a: frame_spi_obj_group_bin_0044 (RW)
0x4b: frame_spi_obj_group_bin_0124 (RW)
0x4c: frame_spi_obj_group_bin_0209 (RW)
0x4d: frame_spi_obj_group_bin_0292 (RW)
0x4e: frame_spi_obj_group_bin_0054 (RW)
0x4f: frame_spi_obj_group_bin_0135 (RW)
0x50: frame_spi_obj_group_bin_0217 (RW)
0x51: frame_spi_obj_group_bin_0301 (RW)
0x52: frame_spi_obj_group_bin_0064 (RW)
0x53: frame_spi_obj_group_bin_0145 (RW)
0x54: frame_spi_obj_group_bin_0227 (RW)
0x55: frame_spi_obj_group_bin_0309 (RW)
0x56: frame_spi_obj_group_bin_0073 (RW)
0x57: frame_spi_obj_group_bin_0155 (RW)
0x58: frame_spi_obj_group_bin_0238 (RW)
0x59: frame_spi_obj_group_bin_0002 (RW)
0x5a: frame_spi_obj_group_bin_0083 (RW)
0x5b: frame_spi_obj_group_bin_0166 (RW)
0x5c: frame_spi_obj_group_bin_0248 (RW)
0x5d: frame_spi_obj_group_bin_0013 (RW)
0x5e: frame_spi_obj_group_bin_0092 (RW)
0x5f: frame_spi_obj_group_bin_0176 (RW)
0x60: frame_spi_obj_group_bin_0258 (RW)
0x61: frame_spi_obj_group_bin_0023 (RW)
0x62: frame_spi_obj_group_bin_0102 (RW)
0x63: frame_spi_obj_group_bin_0186 (RW)
0x64: frame_spi_obj_group_bin_0267 (RW)
0x65: frame_spi_obj_group_bin_0032 (RW)
0x66: frame_spi_obj_group_bin_0113 (RW)
0x67: frame_spi_obj_group_bin_0242 (RW)
0x68: frame_spi_obj_group_bin_0278 (RW)
0x69: frame_spi_obj_group_bin_0041 (RW)
0x6a: frame_spi_obj_group_bin_0122 (RW)
0x6b: frame_spi_obj_group_bin_0207 (RW)
0x6c: frame_spi_obj_group_bin_0290 (RW)
0x6d: frame_spi_obj_group_bin_0051 (RW)
0x6e: frame_spi_obj_group_bin_0132 (RW)
0x6f: frame_spi_obj_group_bin_0215 (RW)
0x70: frame_spi_obj_group_bin_0298 (RW)
0x71: frame_spi_obj_group_bin_0062 (RW)
0x72: frame_spi_obj_group_bin_0141 (RW)
0x73: frame_spi_obj_group_bin_0224 (RW)
0x74: frame_spi_obj_group_bin_0307 (RW)
0x75: frame_spi_obj_group_bin_0071 (RW)
0x76: frame_spi_obj_group_bin_0153 (RW)
0x77: frame_spi_obj_group_bin_0236 (RW)
0x78: frame_spi_obj_group_bin_0316 (RW)
0x79: frame_spi_obj_group_bin_0080 (RW)
0x7a: frame_spi_obj_group_bin_0163 (RW)
0x7b: frame_spi_obj_group_bin_0245 (RW)
0x7c: frame_spi_obj_group_bin_0011 (RW)
0x7d: frame_spi_obj_group_bin_0090 (RW)
0x7e: frame_spi_obj_group_bin_0174 (RW)
0x7f: frame_spi_obj_group_bin_0255 (RW)
0x80: frame_spi_obj_group_bin_0021 (RW)
0x81: frame_spi_obj_group_bin_0100 (RW)
0x82: frame_spi_obj_group_bin_0183 (RW)
0x83: frame_spi_obj_group_bin_0265 (RW)
0x84: frame_spi_obj_group_bin_0029 (RW)
0x85: frame_spi_obj_group_bin_0110 (RW)
0x86: frame_spi_obj_group_bin_0195 (RW)
0x87: frame_spi_obj_group_bin_0275 (RW)
0x88: frame_spi_obj_group_bin_0038 (RW)
0x89: frame_spi_obj_group_bin_0119 (RW)
0x8a: frame_spi_obj_group_bin_0205 (RW)
0x8b: frame_spi_obj_group_bin_0286 (RW)
0x8c: frame_spi_obj_group_bin_0048 (RW)
0x8d: frame_spi_obj_group_bin_0129 (RW)
0x8e: frame_spi_obj_group_bin_0213 (RW)
0x8f: frame_spi_obj_group_bin_0296 (RW)
0x90: frame_spi_obj_group_bin_0060 (RW)
0x91: frame_spi_obj_group_bin_0139 (RW)
0x92: frame_spi_obj_group_bin_0173 (RW)
0x93: frame_spi_obj_group_bin_0264 (RW)
0x94: frame_spi_obj_group_bin_0037 (RW)
0x95: frame_spi_obj_group_bin_0128 (RW)
0x96: frame_spi_obj_group_bin_0221 (RW)
0x97: frame_spi_obj_group_bin_0312 (RW)
0x98: frame_spi_obj_group_bin_0125 (RW)
0x99: frame_spi_obj_group_bin_0268 (RW)
0x9a: frame_spi_obj_group_bin_0243 (RW)
0x9b: frame_spi_obj_group_bin_0046 (RW)
0x9c: frame_spi_obj_group_bin_0137 (RW)
0x9d: frame_spi_obj_group_bin_0201 (RW)
0x9e: frame_spi_obj_group_bin_0024 (RW)
0x9f: frame_spi_obj_group_bin_0164 (RW)
0xa0: frame_spi_obj_group_bin_0190 (RW)
0xa1: frame_spi_obj_group_bin_0281 (RW)
0xa2: frame_spi_obj_group_bin_0055 (RW)
0xa3: frame_spi_obj_group_bin_0146 (RW)
0xa4: frame_spi_obj_group_bin_0107 (RW)
0xa5: frame_spi_obj_group_bin_0192 (RW)
0xa6: frame_spi_obj_group_bin_0273 (RW)
0xa7: frame_spi_obj_group_bin_0036 (RW)
0xa8: frame_spi_obj_group_bin_0117 (RW)
0xa9: frame_spi_obj_group_bin_0203 (RW)
0xaa: frame_spi_obj_group_bin_0283 (RW)
0xab: frame_spi_obj_group_bin_0247 (RW)
0xac: frame_spi_obj_group_bin_0126 (RW)
0xad: frame_spi_obj_group_bin_0211 (RW)
0xae: frame_spi_obj_group_bin_0294 (RW)
0xaf: frame_spi_obj_group_bin_0057 (RW)
0xb0: frame_spi_obj_group_bin_0070 (RW)
0xb1: frame_spi_obj_group_bin_0220 (RW)
0xb2: frame_spi_obj_group_bin_0303 (RW)
0xb3: frame_spi_obj_group_bin_0028 (RW)
0xb4: frame_spi_obj_group_bin_0118 (RW)
0xb5: frame_spi_obj_group_bin_0212 (RW)
0xb6: frame_spi_obj_group_bin_0304 (RW)
0xb7: frame_spi_obj_group_bin_0077 (RW)
0xb8: frame_spi_obj_group_bin_0157 (RW)
0xb9: frame_spi_obj_group_bin_0042 (RW)
0xba: frame_spi_obj_group_bin_0184 (RW)
0xbb: frame_spi_obj_group_bin_0008 (RW)
0xbc: frame_spi_obj_group_bin_0149 (RW)
0xbd: frame_spi_obj_group_bin_0251 (RW)
0xbe: frame_spi_obj_group_bin_0114 (RW)
0xbf: frame_spi_obj_group_bin_0256 (RW)
0xc0: frame_spi_obj_group_bin_0271 (RW)
0xc1: frame_spi_obj_group_bin_0045 (RW)
0xc2: frame_spi_obj_group_bin_0136 (RW)
0xc3: frame_spi_obj_group_bin_0228 (RW)
0xc4: frame_spi_obj_group_bin_0003 (RW)
0xc5: frame_spi_obj_group_bin_0093 (RW)
0xc6: frame_spi_obj_group_bin_0187 (RW)
0xc7: frame_spi_obj_group_bin_0279 (RW)
0xc8: frame_spi_obj_group_bin_0053 (RW)
0xc9: frame_spi_obj_group_bin_0143 (RW)
0xca: frame_spi_obj_group_bin_0237 (RW)
0xcb: frame_spi_obj_group_bin_0012 (RW)
0xcc: frame_spi_obj_group_bin_0101 (RW)
0xcd: frame_spi_obj_group_bin_0197 (RW)
0xce: frame_spi_obj_group_bin_0288 (RW)
0xcf: frame_spi_obj_group_bin_0061 (RW)
0xd0: frame_spi_obj_group_bin_0152 (RW)
0xd1: frame_spi_obj_group_bin_0244 (RW)
0xd2: frame_spi_obj_group_bin_0020 (RW)
0xd3: frame_spi_obj_group_bin_0109 (RW)
0xd4: frame_spi_obj_group_bin_0204 (RW)
0xd5: frame_spi_obj_group_bin_0295 (RW)
0xd6: frame_spi_obj_group_bin_0067 (RW)
0xd7: frame_spi_obj_group_bin_0160 (RW)
0xd8: frame_spi_obj_group_bin_0310 (RW)
0xd9: frame_spi_obj_group_bin_0133 (RW)
0xda: frame_spi_obj_group_bin_0276 (RW)
0xdb: frame_spi_obj_group_bin_0098 (RW)
0xdc: frame_spi_obj_group_bin_0241 (RW)
0xdd: frame_spi_obj_group_bin_0065 (RW)
0xde: frame_spi_obj_group_bin_0208 (RW)
0xdf: frame_spi_obj_group_bin_0030 (RW)
0xe0: frame_spi_obj_group_bin_0035 (RW)
0xe1: frame_spi_obj_group_bin_0314 (RW)
0xe2: frame_spi_obj_group_bin_0218 (RW)
0xe3: frame_spi_obj_group_bin_0282 (RW)
0xe4: frame_spi_obj_group_bin_0084 (RW)
0xe5: frame_spi_obj_group_bin_0177 (RW)
0xe6: frame_spi_obj_group_bin_0069 (RW)
0xe7: frame_spi_obj_group_bin_0198 (RW)
0xe8: frame_spi_obj_group_bin_0134 (RW)
0xe9: frame_spi_obj_group_bin_0226 (RW)
0xea: frame_spi_obj_group_bin_0095 (RW)
0xeb: frame_spi_obj_group_bin_0091 (RW)
0xec: frame_spi_obj_group_bin_0185 (RW)
0xed: frame_spi_obj_group_bin_0277 (RW)
0xee: frame_spi_obj_group_bin_0050 (RW)
0xef: frame_spi_obj_group_bin_0140 (RW)
0xf0: frame_spi_obj_group_bin_0235 (RW)
0xf1: frame_spi_obj_group_bin_0010 (RW)
0xf2: frame_spi_obj_group_bin_0099 (RW)
0xf3: frame_spi_obj_group_bin_0194 (RW)
0xf4: frame_spi_obj_group_bin_0285 (RW)
0xf5: frame_spi_obj_group_bin_0059 (RW)
0xf6: frame_spi_obj_group_bin_0150 (RW)
0xf7: frame_spi_obj_group_bin_0019 (RW)
0xf8: frame_spi_obj_group_bin_0104 (RW)
0xf9: frame_spi_obj_group_bin_0225 (RW)
0xfa: frame_spi_obj_group_bin_0049 (RW)
0xfb: frame_spi_obj_group_bin_0193 (RW)
0xfc: frame_spi_obj_group_bin_0017 (RW)
0xfd: frame_spi_obj_group_bin_0156 (RW)
0xfe: frame_spi_obj_group_bin_0299 (RW)
0xff: frame_spi_obj_group_bin_0120 (RW)
}
pt_spi_obj_group_bin_0247 {
0x0: frame_spi_obj_group_bin_0246 (RW, uncached)
}
pt_timer_obj_group_bin_0000 {
0x100: frame_timer_obj_group_bin_0110 (RW)
0x101: frame_timer_obj_group_bin_0198 (RW)
0x102: frame_timer_obj_group_bin_0286 (RW)
0x103: frame_timer_obj_group_bin_0071 (RW)
0x104: frame_timer_obj_group_bin_0159 (RW)
0x105: frame_timer_obj_group_bin_0246 (RW)
0x106: frame_timer_obj_group_bin_0032 (RW)
0x107: frame_timer_obj_group_bin_0117 (RW)
0x108: frame_timer_obj_group_bin_0204 (RW)
0x109: frame_timer_obj_group_bin_0292 (RW)
0x10: frame_timer_obj_group_bin_0000 (RX)
0x10a: frame_timer_obj_group_bin_0078 (RW)
0x10b: frame_timer_obj_group_bin_0165 (RW)
0x10c: frame_timer_obj_group_bin_0253 (RW)
0x10d: frame_timer_obj_group_bin_0038 (RW)
0x10e: frame_timer_obj_group_bin_0124 (RW)
0x10f: frame_timer_obj_group_bin_0211 (RW)
0x110: frame_timer_obj_group_bin_0299 (RW)
0x111: frame_timer_obj_group_bin_0086 (RW)
0x112: frame_timer_obj_group_bin_0171 (RW)
0x113: frame_timer_obj_group_bin_0260 (RW)
0x114: frame_timer_obj_group_bin_0045 (RW)
0x115: frame_timer_obj_group_bin_0132 (RW)
0x116: frame_timer_obj_group_bin_0219 (RW)
0x117: frame_timer_obj_group_bin_0006 (RW)
0x118: frame_timer_obj_group_bin_0168 (RW)
0x119: frame_timer_obj_group_bin_0160 (RW)
0x11: frame_timer_obj_group_bin_0001 (RX)
0x11a: frame_timer_obj_group_bin_0072 (RW)
0x11b: frame_timer_obj_group_bin_0270 (RW)
0x11c: frame_timer_obj_group_bin_0102 (RW)
0x11d: frame_timer_obj_group_bin_0238 (RW)
0x11e: frame_timer_obj_group_bin_0069 (RW)
0x11f: frame_timer_obj_group_bin_0202 (RW)
0x120: frame_timer_obj_group_bin_0039 (RW)
0x121: frame_timer_obj_group_bin_0059 (RW)
0x122: frame_timer_obj_group_bin_0151 (RW)
0x123: frame_timer_obj_group_bin_0140 (RW)
0x124: frame_timer_obj_group_bin_0237 (RW)
0x125: frame_timer_obj_group_bin_0023 (RW)
0x126: frame_timer_obj_group_bin_0012 (RW)
0x127: frame_timer_obj_group_bin_0050 (RW)
0x128: frame_timer_obj_group_bin_0284 (RW)
0x129: frame_timer_obj_group_bin_0221 (RW)
0x12: frame_timer_obj_group_bin_0210 (RX)
0x12a: frame_timer_obj_group_bin_0157 (RW)
0x12b: frame_timer_obj_group_bin_0244 (RW)
0x12c: frame_timer_obj_group_bin_0030 (RW)
0x12d: frame_timer_obj_group_bin_0115 (RW)
0x12e: frame_timer_obj_group_bin_0207 (RW)
0x12f: frame_timer_obj_group_bin_0290 (RW)
0x131: frame_timer_obj_group_bin_0179 (RW)
0x134: frame_timer_obj_group_bin_0083 (RW)
0x137: frame_timer_obj_group_bin_0084 (RW)
0x13: frame_timer_obj_group_bin_0289 (RX)
0x13a: frame_timer_obj_group_bin_0222 (RW)
0x13b: frame_timer_obj_group_bin_0055 (RW)
0x13c: frame_timer_obj_group_bin_0190 (RW)
0x13d: frame_timer_obj_group_bin_0024 (RW)
0x140: frame_timer_obj_group_bin_0267 (RW)
0x141: frame_timer_obj_group_bin_0053 (RW)
0x142: frame_timer_obj_group_bin_0139 (RW)
0x143: frame_timer_obj_group_bin_0227 (RW)
0x146: frame_timer_obj_group_bin_0187 (RW)
0x147: frame_timer_obj_group_bin_0275 (RW)
0x148: frame_timer_obj_group_bin_0061 (RW)
0x149: frame_timer_obj_group_bin_0147 (RW)
0x14: frame_timer_obj_group_bin_0066 (RX)
0x15: frame_timer_obj_group_bin_0144 (RX)
0x16: frame_timer_obj_group_bin_0220 (RX)
0x17: frame_timer_obj_group_bin_0297 (RX)
0x18: frame_timer_obj_group_bin_0075 (RX)
0x19: frame_timer_obj_group_bin_0079 (RX)
0x1a: frame_timer_obj_group_bin_0155 (RX)
0x1b: frame_timer_obj_group_bin_0007 (RX)
0x1c: frame_timer_obj_group_bin_0085 (RX)
0x1d: frame_timer_obj_group_bin_0162 (RX)
0x2d: frame_timer_obj_group_bin_0199 (RW)
0x2e: frame_timer_obj_group_bin_0278 (RW)
0x2f: frame_timer_obj_group_bin_0054 (RW)
0x30: frame_timer_obj_group_bin_0004 (RW)
0x31: frame_timer_obj_group_bin_0208 (RW)
0x32: frame_timer_obj_group_bin_0287 (RW)
0x33: frame_timer_obj_group_bin_0064 (RW)
0x34: frame_timer_obj_group_bin_0141 (RW)
0x35: frame_timer_obj_group_bin_0217 (RW)
0x36: frame_timer_obj_group_bin_0295 (RW)
0x37: frame_timer_obj_group_bin_0073 (RW)
0x38: frame_timer_obj_group_bin_0150 (RW)
0x39: frame_timer_obj_group_bin_0228 (RW)
0x3a: frame_timer_obj_group_bin_0005 (RW)
0x3b: frame_timer_obj_group_bin_0082 (RW)
0x3c: frame_timer_obj_group_bin_0161 (RW)
0x3d: frame_timer_obj_group_bin_0239 (RW)
0x3e: frame_timer_obj_group_bin_0016 (RW)
0x3f: frame_timer_obj_group_bin_0091 (RW)
0x40: frame_timer_obj_group_bin_0169 (RW)
0x41: frame_timer_obj_group_bin_0248 (RW)
0x42: frame_timer_obj_group_bin_0025 (RW)
0x43: frame_timer_obj_group_bin_0101 (RW)
0x44: frame_timer_obj_group_bin_0178 (RW)
0x45: frame_timer_obj_group_bin_0257 (RW)
0x46: frame_timer_obj_group_bin_0033 (RW)
0x47: frame_timer_obj_group_bin_0109 (RW)
0x48: frame_timer_obj_group_bin_0188 (RW)
0x49: frame_timer_obj_group_bin_0266 (RW)
0x4a: frame_timer_obj_group_bin_0042 (RW)
0x4b: frame_timer_obj_group_bin_0118 (RW)
0x4c: frame_timer_obj_group_bin_0197 (RW)
0x4d: frame_timer_obj_group_bin_0276 (RW)
0x4e: frame_timer_obj_group_bin_0052 (RW)
0x4f: frame_timer_obj_group_bin_0128 (RW)
0x50: frame_timer_obj_group_bin_0205 (RW)
0x51: frame_timer_obj_group_bin_0285 (RW)
0x52: frame_timer_obj_group_bin_0062 (RW)
0x53: frame_timer_obj_group_bin_0138 (RW)
0x54: frame_timer_obj_group_bin_0215 (RW)
0x55: frame_timer_obj_group_bin_0293 (RW)
0x56: frame_timer_obj_group_bin_0070 (RW)
0x57: frame_timer_obj_group_bin_0148 (RW)
0x58: frame_timer_obj_group_bin_0226 (RW)
0x59: frame_timer_obj_group_bin_0002 (RW)
0x5a: frame_timer_obj_group_bin_0080 (RW)
0x5b: frame_timer_obj_group_bin_0158 (RW)
0x5c: frame_timer_obj_group_bin_0236 (RW)
0x5d: frame_timer_obj_group_bin_0014 (RW)
0x5e: frame_timer_obj_group_bin_0089 (RW)
0x5f: frame_timer_obj_group_bin_0166 (RW)
0x60: frame_timer_obj_group_bin_0245 (RW)
0x61: frame_timer_obj_group_bin_0022 (RW)
0x62: frame_timer_obj_group_bin_0098 (RW)
0x63: frame_timer_obj_group_bin_0175 (RW)
0x64: frame_timer_obj_group_bin_0254 (RW)
0x65: frame_timer_obj_group_bin_0031 (RW)
0x66: frame_timer_obj_group_bin_0107 (RW)
0x67: frame_timer_obj_group_bin_0230 (RW)
0x68: frame_timer_obj_group_bin_0264 (RW)
0x69: frame_timer_obj_group_bin_0040 (RW)
0x6a: frame_timer_obj_group_bin_0116 (RW)
0x6b: frame_timer_obj_group_bin_0195 (RW)
0x6c: frame_timer_obj_group_bin_0274 (RW)
0x6d: frame_timer_obj_group_bin_0049 (RW)
0x6e: frame_timer_obj_group_bin_0125 (RW)
0x6f: frame_timer_obj_group_bin_0203 (RW)
0x70: frame_timer_obj_group_bin_0282 (RW)
0x71: frame_timer_obj_group_bin_0060 (RW)
0x72: frame_timer_obj_group_bin_0135 (RW)
0x73: frame_timer_obj_group_bin_0212 (RW)
0x74: frame_timer_obj_group_bin_0291 (RW)
0x75: frame_timer_obj_group_bin_0068 (RW)
0x76: frame_timer_obj_group_bin_0146 (RW)
0x77: frame_timer_obj_group_bin_0224 (RW)
0x78: frame_timer_obj_group_bin_0300 (RW)
0x79: frame_timer_obj_group_bin_0077 (RW)
0x7a: frame_timer_obj_group_bin_0156 (RW)
0x7b: frame_timer_obj_group_bin_0233 (RW)
0x7c: frame_timer_obj_group_bin_0011 (RW)
0x7d: frame_timer_obj_group_bin_0087 (RW)
0x7e: frame_timer_obj_group_bin_0164 (RW)
0x7f: frame_timer_obj_group_bin_0242 (RW)
0x80: frame_timer_obj_group_bin_0021 (RW)
0x81: frame_timer_obj_group_bin_0096 (RW)
0x82: frame_timer_obj_group_bin_0172 (RW)
0x83: frame_timer_obj_group_bin_0252 (RW)
0x84: frame_timer_obj_group_bin_0028 (RW)
0x85: frame_timer_obj_group_bin_0105 (RW)
0x86: frame_timer_obj_group_bin_0183 (RW)
0x87: frame_timer_obj_group_bin_0261 (RW)
0x88: frame_timer_obj_group_bin_0037 (RW)
0x89: frame_timer_obj_group_bin_0113 (RW)
0x8a: frame_timer_obj_group_bin_0193 (RW)
0x8b: frame_timer_obj_group_bin_0272 (RW)
0x8c: frame_timer_obj_group_bin_0046 (RW)
0x8d: frame_timer_obj_group_bin_0123 (RW)
0x8e: frame_timer_obj_group_bin_0201 (RW)
0x8f: frame_timer_obj_group_bin_0280 (RW)
0x90: frame_timer_obj_group_bin_0057 (RW)
0x91: frame_timer_obj_group_bin_0133 (RW)
0x92: frame_timer_obj_group_bin_0163 (RW)
0x93: frame_timer_obj_group_bin_0251 (RW)
0x94: frame_timer_obj_group_bin_0036 (RW)
0x95: frame_timer_obj_group_bin_0122 (RW)
0x96: frame_timer_obj_group_bin_0209 (RW)
0x97: frame_timer_obj_group_bin_0296 (RW)
0x98: frame_timer_obj_group_bin_0119 (RW)
0x99: frame_timer_obj_group_bin_0154 (RW)
0x9a: frame_timer_obj_group_bin_0231 (RW)
0x9b: frame_timer_obj_group_bin_0044 (RW)
0x9c: frame_timer_obj_group_bin_0130 (RW)
0x9d: frame_timer_obj_group_bin_0189 (RW)
0x9e: frame_timer_obj_group_bin_0240 (RW)
0x9f: frame_timer_obj_group_bin_0018 (RW)
0xa0: frame_timer_obj_group_bin_0093 (RW)
0xa1: frame_timer_obj_group_bin_0170 (RW)
0xa2: frame_timer_obj_group_bin_0250 (RW)
0xa3: frame_timer_obj_group_bin_0026 (RW)
0xa4: frame_timer_obj_group_bin_0103 (RW)
0xa5: frame_timer_obj_group_bin_0180 (RW)
0xa6: frame_timer_obj_group_bin_0259 (RW)
0xa7: frame_timer_obj_group_bin_0035 (RW)
0xa8: frame_timer_obj_group_bin_0111 (RW)
0xa9: frame_timer_obj_group_bin_0191 (RW)
0xaa: frame_timer_obj_group_bin_0269 (RW)
0xab: frame_timer_obj_group_bin_0235 (RW)
0xac: frame_timer_obj_group_bin_0120 (RW)
0xad: frame_timer_obj_group_bin_0106 (RW)
0xae: frame_timer_obj_group_bin_0194 (RW)
0xaf: frame_timer_obj_group_bin_0281 (RW)
0xb0: frame_timer_obj_group_bin_0067 (RW)
0xb1: frame_timer_obj_group_bin_0243 (RW)
0xb2: frame_timer_obj_group_bin_0241 (RW)
0xb3: frame_timer_obj_group_bin_0027 (RW)
0xb4: frame_timer_obj_group_bin_0112 (RW)
0xb5: frame_timer_obj_group_bin_0200 (RW)
0xb6: frame_timer_obj_group_bin_0288 (RW)
0xb7: frame_timer_obj_group_bin_0074 (RW)
0xb8: frame_timer_obj_group_bin_0206 (RW)
0xb9: frame_timer_obj_group_bin_0041 (RW)
0xba: frame_timer_obj_group_bin_0173 (RW)
0xbb: frame_timer_obj_group_bin_0008 (RW)
0xbc: frame_timer_obj_group_bin_0142 (RW)
0xbd: frame_timer_obj_group_bin_0277 (RW)
0xbe: frame_timer_obj_group_bin_0108 (RW)
0xbf: frame_timer_obj_group_bin_0009 (RW)
0xc0: frame_timer_obj_group_bin_0258 (RW)
0xc1: frame_timer_obj_group_bin_0043 (RW)
0xc2: frame_timer_obj_group_bin_0129 (RW)
0xc3: frame_timer_obj_group_bin_0216 (RW)
0xc4: frame_timer_obj_group_bin_0003 (RW)
0xc5: frame_timer_obj_group_bin_0090 (RW)
0xc6: frame_timer_obj_group_bin_0176 (RW)
0xc7: frame_timer_obj_group_bin_0265 (RW)
0xc8: frame_timer_obj_group_bin_0051 (RW)
0xc9: frame_timer_obj_group_bin_0136 (RW)
0xca: frame_timer_obj_group_bin_0225 (RW)
0xcb: frame_timer_obj_group_bin_0013 (RW)
0xcc: frame_timer_obj_group_bin_0097 (RW)
0xcd: frame_timer_obj_group_bin_0185 (RW)
0xce: frame_timer_obj_group_bin_0273 (RW)
0xcf: frame_timer_obj_group_bin_0058 (RW)
0xd0: frame_timer_obj_group_bin_0145 (RW)
0xd1: frame_timer_obj_group_bin_0232 (RW)
0xd2: frame_timer_obj_group_bin_0020 (RW)
0xd3: frame_timer_obj_group_bin_0104 (RW)
0xd4: frame_timer_obj_group_bin_0192 (RW)
0xd5: frame_timer_obj_group_bin_0279 (RW)
0xd6: frame_timer_obj_group_bin_0065 (RW)
0xd7: frame_timer_obj_group_bin_0153 (RW)
0xd8: frame_timer_obj_group_bin_0294 (RW)
0xd9: frame_timer_obj_group_bin_0126 (RW)
0xda: frame_timer_obj_group_bin_0262 (RW)
0xdb: frame_timer_obj_group_bin_0094 (RW)
0xdc: frame_timer_obj_group_bin_0229 (RW)
0xdd: frame_timer_obj_group_bin_0063 (RW)
0xde: frame_timer_obj_group_bin_0196 (RW)
0xdf: frame_timer_obj_group_bin_0029 (RW)
0xe0: frame_timer_obj_group_bin_0034 (RW)
0xe1: frame_timer_obj_group_bin_0298 (RW)
0xe2: frame_timer_obj_group_bin_0131 (RW)
0xe3: frame_timer_obj_group_bin_0268 (RW)
0xe4: frame_timer_obj_group_bin_0081 (RW)
0xe5: frame_timer_obj_group_bin_0167 (RW)
0xe6: frame_timer_obj_group_bin_0255 (RW)
0xe7: frame_timer_obj_group_bin_0186 (RW)
0xe8: frame_timer_obj_group_bin_0127 (RW)
0xe9: frame_timer_obj_group_bin_0214 (RW)
0xea: frame_timer_obj_group_bin_0092 (RW)
0xeb: frame_timer_obj_group_bin_0088 (RW)
0xec: frame_timer_obj_group_bin_0174 (RW)
0xed: frame_timer_obj_group_bin_0263 (RW)
0xee: frame_timer_obj_group_bin_0048 (RW)
0xef: frame_timer_obj_group_bin_0134 (RW)
0xf0: frame_timer_obj_group_bin_0223 (RW)
0xf1: frame_timer_obj_group_bin_0010 (RW)
0xf2: frame_timer_obj_group_bin_0095 (RW)
0xf3: frame_timer_obj_group_bin_0182 (RW)
0xf4: frame_timer_obj_group_bin_0271 (RW)
0xf5: frame_timer_obj_group_bin_0056 (RW)
0xf6: frame_timer_obj_group_bin_0143 (RW)
0xf7: frame_timer_obj_group_bin_0019 (RW)
0xf8: frame_timer_obj_group_bin_0100 (RW)
0xf9: frame_timer_obj_group_bin_0213 (RW)
0xfa: frame_timer_obj_group_bin_0047 (RW)
0xfb: frame_timer_obj_group_bin_0181 (RW)
0xfc: frame_timer_obj_group_bin_0017 (RW)
0xfd: frame_timer_obj_group_bin_0149 (RW)
0xfe: frame_timer_obj_group_bin_0283 (RW)
0xff: frame_timer_obj_group_bin_0114 (RW)
}
pt_timer_obj_group_bin_0235 {
0x0: frame_timer_obj_group_bin_0234 (RW, uncached)
}
pt_uart_gcs_group_bin_0000 {
0x100: frame_uart_gcs_group_bin_0116 (RW)
0x101: frame_uart_gcs_group_bin_0209 (RW)
0x102: frame_uart_gcs_group_bin_0299 (RW)
0x103: frame_uart_gcs_group_bin_0075 (RW)
0x104: frame_uart_gcs_group_bin_0167 (RW)
0x105: frame_uart_gcs_group_bin_0258 (RW)
0x106: frame_uart_gcs_group_bin_0034 (RW)
0x107: frame_uart_gcs_group_bin_0123 (RW)
0x108: frame_uart_gcs_group_bin_0215 (RW)
0x109: frame_uart_gcs_group_bin_0305 (RW)
0x10: frame_uart_gcs_group_bin_0000 (RX)
0x10a: frame_uart_gcs_group_bin_0082 (RW)
0x10b: frame_uart_gcs_group_bin_0174 (RW)
0x10c: frame_uart_gcs_group_bin_0265 (RW)
0x10d: frame_uart_gcs_group_bin_0040 (RW)
0x10e: frame_uart_gcs_group_bin_0130 (RW)
0x10f: frame_uart_gcs_group_bin_0222 (RW)
0x110: frame_uart_gcs_group_bin_0312 (RW)
0x111: frame_uart_gcs_group_bin_0090 (RW)
0x112: frame_uart_gcs_group_bin_0181 (RW)
0x113: frame_uart_gcs_group_bin_0272 (RW)
0x114: frame_uart_gcs_group_bin_0047 (RW)
0x115: frame_uart_gcs_group_bin_0138 (RW)
0x116: frame_uart_gcs_group_bin_0230 (RW)
0x117: frame_uart_gcs_group_bin_0006 (RW)
0x118: frame_uart_gcs_group_bin_0177 (RW)
0x119: frame_uart_gcs_group_bin_0168 (RW)
0x11: frame_uart_gcs_group_bin_0001 (RX)
0x11a: frame_uart_gcs_group_bin_0076 (RW)
0x11b: frame_uart_gcs_group_bin_0282 (RW)
0x11c: frame_uart_gcs_group_bin_0106 (RW)
0x11d: frame_uart_gcs_group_bin_0249 (RW)
0x11e: frame_uart_gcs_group_bin_0073 (RW)
0x11f: frame_uart_gcs_group_bin_0213 (RW)
0x120: frame_uart_gcs_group_bin_0041 (RW)
0x121: frame_uart_gcs_group_bin_0062 (RW)
0x122: frame_uart_gcs_group_bin_0158 (RW)
0x123: frame_uart_gcs_group_bin_0147 (RW)
0x124: frame_uart_gcs_group_bin_0248 (RW)
0x125: frame_uart_gcs_group_bin_0112 (RW)
0x126: frame_uart_gcs_group_bin_0012 (RW)
0x127: frame_uart_gcs_group_bin_0052 (RW)
0x128: frame_uart_gcs_group_bin_0297 (RW)
0x129: frame_uart_gcs_group_bin_0232 (RW)
0x12: frame_uart_gcs_group_bin_0221 (RX)
0x12a: frame_uart_gcs_group_bin_0165 (RW)
0x12b: frame_uart_gcs_group_bin_0256 (RW)
0x12c: frame_uart_gcs_group_bin_0032 (RW)
0x12d: frame_uart_gcs_group_bin_0121 (RW)
0x12e: frame_uart_gcs_group_bin_0218 (RW)
0x12f: frame_uart_gcs_group_bin_0303 (RW)
0x130: frame_uart_gcs_group_bin_0080 (RW)
0x131: frame_uart_gcs_group_bin_0190 (RW)
0x132: frame_uart_gcs_group_bin_0261 (RW)
0x134: frame_uart_gcs_group_bin_0087 (RW)
0x137: frame_uart_gcs_group_bin_0088 (RW)
0x13: frame_uart_gcs_group_bin_0302 (RX)
0x13a: frame_uart_gcs_group_bin_0233 (RW)
0x13d: frame_uart_gcs_group_bin_0026 (RW)
0x140: frame_uart_gcs_group_bin_0279 (RW)
0x141: frame_uart_gcs_group_bin_0055 (RW)
0x142: frame_uart_gcs_group_bin_0146 (RW)
0x143: frame_uart_gcs_group_bin_0238 (RW)
0x146: frame_uart_gcs_group_bin_0198 (RW)
0x147: frame_uart_gcs_group_bin_0288 (RW)
0x148: frame_uart_gcs_group_bin_0064 (RW)
0x149: frame_uart_gcs_group_bin_0154 (RW)
0x14: frame_uart_gcs_group_bin_0069 (RX)
0x14c: frame_uart_gcs_group_bin_0111 (RW)
0x14d: frame_uart_gcs_group_bin_0205 (RW)
0x14e: frame_uart_gcs_group_bin_0294 (RW)
0x14f: frame_uart_gcs_group_bin_0070 (RW)
0x152: frame_uart_gcs_group_bin_0142 (RW)
0x153: frame_uart_gcs_group_bin_0285 (RW)
0x154: frame_uart_gcs_group_bin_0108 (RW)
0x155: frame_uart_gcs_group_bin_0251 (RW)
0x157: frame_uart_gcs_group_bin_0170 (RWX)
0x15: frame_uart_gcs_group_bin_0151 (RX)
0x16: frame_uart_gcs_group_bin_0231 (RX)
0x17: frame_uart_gcs_group_bin_0310 (RX)
0x18: frame_uart_gcs_group_bin_0079 (RX)
0x19: frame_uart_gcs_group_bin_0083 (RX)
0x1a: frame_uart_gcs_group_bin_0162 (RX)
0x1b: frame_uart_gcs_group_bin_0007 (RX)
0x1c: frame_uart_gcs_group_bin_0089 (RX)
0x1d: frame_uart_gcs_group_bin_0171 (RX)
0x1e: frame_uart_gcs_group_bin_0252 (RX)
0x1f: frame_uart_gcs_group_bin_0019 (RX)
0x20: frame_uart_gcs_group_bin_0097 (RX)
0x30: frame_uart_gcs_group_bin_0004 (RW)
0x31: frame_uart_gcs_group_bin_0219 (RW)
0x32: frame_uart_gcs_group_bin_0300 (RW)
0x33: frame_uart_gcs_group_bin_0067 (RW)
0x34: frame_uart_gcs_group_bin_0148 (RW)
0x35: frame_uart_gcs_group_bin_0228 (RW)
0x36: frame_uart_gcs_group_bin_0308 (RW)
0x37: frame_uart_gcs_group_bin_0077 (RW)
0x38: frame_uart_gcs_group_bin_0157 (RW)
0x39: frame_uart_gcs_group_bin_0239 (RW)
0x3a: frame_uart_gcs_group_bin_0005 (RW)
0x3b: frame_uart_gcs_group_bin_0086 (RW)
0x3c: frame_uart_gcs_group_bin_0169 (RW)
0x3d: frame_uart_gcs_group_bin_0250 (RW)
0x3e: frame_uart_gcs_group_bin_0017 (RW)
0x3f: frame_uart_gcs_group_bin_0095 (RW)
0x40: frame_uart_gcs_group_bin_0178 (RW)
0x41: frame_uart_gcs_group_bin_0260 (RW)
0x42: frame_uart_gcs_group_bin_0027 (RW)
0x43: frame_uart_gcs_group_bin_0105 (RW)
0x44: frame_uart_gcs_group_bin_0188 (RW)
0x45: frame_uart_gcs_group_bin_0269 (RW)
0x46: frame_uart_gcs_group_bin_0035 (RW)
0x47: frame_uart_gcs_group_bin_0115 (RW)
0x48: frame_uart_gcs_group_bin_0199 (RW)
0x49: frame_uart_gcs_group_bin_0278 (RW)
0x4a: frame_uart_gcs_group_bin_0044 (RW)
0x4b: frame_uart_gcs_group_bin_0124 (RW)
0x4c: frame_uart_gcs_group_bin_0208 (RW)
0x4d: frame_uart_gcs_group_bin_0289 (RW)
0x4e: frame_uart_gcs_group_bin_0054 (RW)
0x4f: frame_uart_gcs_group_bin_0134 (RW)
0x50: frame_uart_gcs_group_bin_0216 (RW)
0x51: frame_uart_gcs_group_bin_0298 (RW)
0x52: frame_uart_gcs_group_bin_0065 (RW)
0x53: frame_uart_gcs_group_bin_0145 (RW)
0x54: frame_uart_gcs_group_bin_0226 (RW)
0x55: frame_uart_gcs_group_bin_0306 (RW)
0x56: frame_uart_gcs_group_bin_0074 (RW)
0x57: frame_uart_gcs_group_bin_0155 (RW)
0x58: frame_uart_gcs_group_bin_0237 (RW)
0x59: frame_uart_gcs_group_bin_0002 (RW)
0x5a: frame_uart_gcs_group_bin_0084 (RW)
0x5b: frame_uart_gcs_group_bin_0166 (RW)
0x5c: frame_uart_gcs_group_bin_0247 (RW)
0x5d: frame_uart_gcs_group_bin_0014 (RW)
0x5e: frame_uart_gcs_group_bin_0093 (RW)
0x5f: frame_uart_gcs_group_bin_0175 (RW)
0x60: frame_uart_gcs_group_bin_0257 (RW)
0x61: frame_uart_gcs_group_bin_0024 (RW)
0x62: frame_uart_gcs_group_bin_0102 (RW)
0x63: frame_uart_gcs_group_bin_0185 (RW)
0x64: frame_uart_gcs_group_bin_0266 (RW)
0x65: frame_uart_gcs_group_bin_0033 (RW)
0x66: frame_uart_gcs_group_bin_0113 (RW)
0x67: frame_uart_gcs_group_bin_0241 (RW)
0x68: frame_uart_gcs_group_bin_0276 (RW)
0x69: frame_uart_gcs_group_bin_0042 (RW)
0x6a: frame_uart_gcs_group_bin_0122 (RW)
0x6b: frame_uart_gcs_group_bin_0206 (RW)
0x6c: frame_uart_gcs_group_bin_0287 (RW)
0x6d: frame_uart_gcs_group_bin_0051 (RW)
0x6e: frame_uart_gcs_group_bin_0131 (RW)
0x6f: frame_uart_gcs_group_bin_0214 (RW)
0x70: frame_uart_gcs_group_bin_0295 (RW)
0x71: frame_uart_gcs_group_bin_0063 (RW)
0x72: frame_uart_gcs_group_bin_0141 (RW)
0x73: frame_uart_gcs_group_bin_0223 (RW)
0x74: frame_uart_gcs_group_bin_0304 (RW)
0x75: frame_uart_gcs_group_bin_0072 (RW)
0x76: frame_uart_gcs_group_bin_0153 (RW)
0x77: frame_uart_gcs_group_bin_0235 (RW)
0x78: frame_uart_gcs_group_bin_0313 (RW)
0x79: frame_uart_gcs_group_bin_0081 (RW)
0x7a: frame_uart_gcs_group_bin_0163 (RW)
0x7b: frame_uart_gcs_group_bin_0244 (RW)
0x7c: frame_uart_gcs_group_bin_0011 (RW)
0x7d: frame_uart_gcs_group_bin_0091 (RW)
0x7e: frame_uart_gcs_group_bin_0173 (RW)
0x7f: frame_uart_gcs_group_bin_0254 (RW)
0x80: frame_uart_gcs_group_bin_0022 (RW)
0x81: frame_uart_gcs_group_bin_0100 (RW)
0x82: frame_uart_gcs_group_bin_0182 (RW)
0x83: frame_uart_gcs_group_bin_0264 (RW)
0x84: frame_uart_gcs_group_bin_0030 (RW)
0x85: frame_uart_gcs_group_bin_0110 (RW)
0x86: frame_uart_gcs_group_bin_0194 (RW)
0x87: frame_uart_gcs_group_bin_0273 (RW)
0x88: frame_uart_gcs_group_bin_0039 (RW)
0x89: frame_uart_gcs_group_bin_0119 (RW)
0x8a: frame_uart_gcs_group_bin_0204 (RW)
0x8b: frame_uart_gcs_group_bin_0284 (RW)
0x8c: frame_uart_gcs_group_bin_0048 (RW)
0x8d: frame_uart_gcs_group_bin_0129 (RW)
0x8e: frame_uart_gcs_group_bin_0212 (RW)
0x8f: frame_uart_gcs_group_bin_0293 (RW)
0x90: frame_uart_gcs_group_bin_0060 (RW)
0x91: frame_uart_gcs_group_bin_0139 (RW)
0x92: frame_uart_gcs_group_bin_0172 (RW)
0x93: frame_uart_gcs_group_bin_0263 (RW)
0x94: frame_uart_gcs_group_bin_0038 (RW)
0x95: frame_uart_gcs_group_bin_0128 (RW)
0x96: frame_uart_gcs_group_bin_0220 (RW)
0x97: frame_uart_gcs_group_bin_0309 (RW)
0x98: frame_uart_gcs_group_bin_0125 (RW)
0x99: frame_uart_gcs_group_bin_0161 (RW)
0x9a: frame_uart_gcs_group_bin_0242 (RW)
0x9b: frame_uart_gcs_group_bin_0046 (RW)
0x9c: frame_uart_gcs_group_bin_0136 (RW)
0x9d: frame_uart_gcs_group_bin_0200 (RW)
0x9e: frame_uart_gcs_group_bin_0025 (RW)
0x9f: frame_uart_gcs_group_bin_0164 (RW)
0xa0: frame_uart_gcs_group_bin_0189 (RW)
0xa1: frame_uart_gcs_group_bin_0180 (RW)
0xa2: frame_uart_gcs_group_bin_0262 (RW)
0xa3: frame_uart_gcs_group_bin_0028 (RW)
0xa4: frame_uart_gcs_group_bin_0107 (RW)
0xa5: frame_uart_gcs_group_bin_0191 (RW)
0xa6: frame_uart_gcs_group_bin_0271 (RW)
0xa7: frame_uart_gcs_group_bin_0037 (RW)
0xa8: frame_uart_gcs_group_bin_0117 (RW)
0xa9: frame_uart_gcs_group_bin_0202 (RW)
0xaa: frame_uart_gcs_group_bin_0281 (RW)
0xab: frame_uart_gcs_group_bin_0246 (RW)
0xac: frame_uart_gcs_group_bin_0126 (RW)
0xad: frame_uart_gcs_group_bin_0210 (RW)
0xae: frame_uart_gcs_group_bin_0291 (RW)
0xaf: frame_uart_gcs_group_bin_0057 (RW)
0xb0: frame_uart_gcs_group_bin_0071 (RW)
0xb1: frame_uart_gcs_group_bin_0255 (RW)
0xb2: frame_uart_gcs_group_bin_0253 (RW)
0xb3: frame_uart_gcs_group_bin_0029 (RW)
0xb4: frame_uart_gcs_group_bin_0118 (RW)
0xb5: frame_uart_gcs_group_bin_0211 (RW)
0xb6: frame_uart_gcs_group_bin_0301 (RW)
0xb7: frame_uart_gcs_group_bin_0078 (RW)
0xb8: frame_uart_gcs_group_bin_0217 (RW)
0xb9: frame_uart_gcs_group_bin_0043 (RW)
0xba: frame_uart_gcs_group_bin_0183 (RW)
0xbb: frame_uart_gcs_group_bin_0008 (RW)
0xbc: frame_uart_gcs_group_bin_0149 (RW)
0xbd: frame_uart_gcs_group_bin_0290 (RW)
0xbe: frame_uart_gcs_group_bin_0114 (RW)
0xbf: frame_uart_gcs_group_bin_0009 (RW)
0xc0: frame_uart_gcs_group_bin_0270 (RW)
0xc1: frame_uart_gcs_group_bin_0045 (RW)
0xc2: frame_uart_gcs_group_bin_0135 (RW)
0xc3: frame_uart_gcs_group_bin_0227 (RW)
0xc4: frame_uart_gcs_group_bin_0003 (RW)
0xc5: frame_uart_gcs_group_bin_0094 (RW)
0xc6: frame_uart_gcs_group_bin_0186 (RW)
0xc7: frame_uart_gcs_group_bin_0277 (RW)
0xc8: frame_uart_gcs_group_bin_0053 (RW)
0xc9: frame_uart_gcs_group_bin_0143 (RW)
0xca: frame_uart_gcs_group_bin_0236 (RW)
0xcb: frame_uart_gcs_group_bin_0013 (RW)
0xcc: frame_uart_gcs_group_bin_0101 (RW)
0xcd: frame_uart_gcs_group_bin_0196 (RW)
0xce: frame_uart_gcs_group_bin_0286 (RW)
0xcf: frame_uart_gcs_group_bin_0061 (RW)
0xd0: frame_uart_gcs_group_bin_0152 (RW)
0xd1: frame_uart_gcs_group_bin_0243 (RW)
0xd2: frame_uart_gcs_group_bin_0021 (RW)
0xd3: frame_uart_gcs_group_bin_0109 (RW)
0xd4: frame_uart_gcs_group_bin_0203 (RW)
0xd5: frame_uart_gcs_group_bin_0292 (RW)
0xd6: frame_uart_gcs_group_bin_0068 (RW)
0xd7: frame_uart_gcs_group_bin_0160 (RW)
0xd8: frame_uart_gcs_group_bin_0307 (RW)
0xd9: frame_uart_gcs_group_bin_0132 (RW)
0xda: frame_uart_gcs_group_bin_0274 (RW)
0xdb: frame_uart_gcs_group_bin_0098 (RW)
0xdc: frame_uart_gcs_group_bin_0240 (RW)
0xdd: frame_uart_gcs_group_bin_0066 (RW)
0xde: frame_uart_gcs_group_bin_0207 (RW)
0xdf: frame_uart_gcs_group_bin_0031 (RW)
0xe0: frame_uart_gcs_group_bin_0036 (RW)
0xe1: frame_uart_gcs_group_bin_0311 (RW)
0xe2: frame_uart_gcs_group_bin_0137 (RW)
0xe3: frame_uart_gcs_group_bin_0280 (RW)
0xe4: frame_uart_gcs_group_bin_0085 (RW)
0xe5: frame_uart_gcs_group_bin_0176 (RW)
0xe6: frame_uart_gcs_group_bin_0267 (RW)
0xe7: frame_uart_gcs_group_bin_0197 (RW)
0xe8: frame_uart_gcs_group_bin_0133 (RW)
0xe9: frame_uart_gcs_group_bin_0225 (RW)
0xea: frame_uart_gcs_group_bin_0096 (RW)
0xeb: frame_uart_gcs_group_bin_0092 (RW)
0xec: frame_uart_gcs_group_bin_0184 (RW)
0xed: frame_uart_gcs_group_bin_0275 (RW)
0xee: frame_uart_gcs_group_bin_0050 (RW)
0xef: frame_uart_gcs_group_bin_0140 (RW)
0xf0: frame_uart_gcs_group_bin_0234 (RW)
0xf1: frame_uart_gcs_group_bin_0010 (RW)
0xf2: frame_uart_gcs_group_bin_0099 (RW)
0xf3: frame_uart_gcs_group_bin_0193 (RW)
0xf4: frame_uart_gcs_group_bin_0283 (RW)
0xf5: frame_uart_gcs_group_bin_0059 (RW)
0xf6: frame_uart_gcs_group_bin_0150 (RW)
0xf7: frame_uart_gcs_group_bin_0020 (RW)
0xf8: frame_uart_gcs_group_bin_0104 (RW)
0xf9: frame_uart_gcs_group_bin_0224 (RW)
0xfa: frame_uart_gcs_group_bin_0049 (RW)
0xfb: frame_uart_gcs_group_bin_0192 (RW)
0xfc: frame_uart_gcs_group_bin_0018 (RW)
0xfd: frame_uart_gcs_group_bin_0156 (RW)
0xfe: frame_uart_gcs_group_bin_0296 (RW)
0xff: frame_uart_gcs_group_bin_0120 (RW)
}
pt_uart_gcs_group_bin_0246 {
0x0: frame_uart_gcs_group_bin_0245 (RW, uncached)
}
pt_uart_px4_group_bin_0000 {
0x100: frame_uart_px4_group_bin_0116 (RW)
0x101: frame_uart_px4_group_bin_0209 (RW)
0x102: frame_uart_px4_group_bin_0299 (RW)
0x103: frame_uart_px4_group_bin_0075 (RW)
0x104: frame_uart_px4_group_bin_0167 (RW)
0x105: frame_uart_px4_group_bin_0258 (RW)
0x106: frame_uart_px4_group_bin_0034 (RW)
0x107: frame_uart_px4_group_bin_0123 (RW)
0x108: frame_uart_px4_group_bin_0215 (RW)
0x109: frame_uart_px4_group_bin_0305 (RW)
0x10: frame_uart_px4_group_bin_0000 (RX)
0x10a: frame_uart_px4_group_bin_0082 (RW)
0x10b: frame_uart_px4_group_bin_0174 (RW)
0x10c: frame_uart_px4_group_bin_0265 (RW)
0x10d: frame_uart_px4_group_bin_0040 (RW)
0x10e: frame_uart_px4_group_bin_0130 (RW)
0x10f: frame_uart_px4_group_bin_0222 (RW)
0x110: frame_uart_px4_group_bin_0312 (RW)
0x111: frame_uart_px4_group_bin_0090 (RW)
0x112: frame_uart_px4_group_bin_0181 (RW)
0x113: frame_uart_px4_group_bin_0272 (RW)
0x114: frame_uart_px4_group_bin_0047 (RW)
0x115: frame_uart_px4_group_bin_0138 (RW)
0x116: frame_uart_px4_group_bin_0230 (RW)
0x117: frame_uart_px4_group_bin_0006 (RW)
0x118: frame_uart_px4_group_bin_0177 (RW)
0x119: frame_uart_px4_group_bin_0168 (RW)
0x11: frame_uart_px4_group_bin_0001 (RX)
0x11a: frame_uart_px4_group_bin_0076 (RW)
0x11b: frame_uart_px4_group_bin_0282 (RW)
0x11c: frame_uart_px4_group_bin_0106 (RW)
0x11d: frame_uart_px4_group_bin_0249 (RW)
0x11e: frame_uart_px4_group_bin_0073 (RW)
0x11f: frame_uart_px4_group_bin_0213 (RW)
0x120: frame_uart_px4_group_bin_0041 (RW)
0x121: frame_uart_px4_group_bin_0062 (RW)
0x122: frame_uart_px4_group_bin_0158 (RW)
0x123: frame_uart_px4_group_bin_0147 (RW)
0x124: frame_uart_px4_group_bin_0248 (RW)
0x125: frame_uart_px4_group_bin_0112 (RW)
0x126: frame_uart_px4_group_bin_0012 (RW)
0x127: frame_uart_px4_group_bin_0052 (RW)
0x128: frame_uart_px4_group_bin_0297 (RW)
0x129: frame_uart_px4_group_bin_0232 (RW)
0x12: frame_uart_px4_group_bin_0221 (RX)
0x12a: frame_uart_px4_group_bin_0165 (RW)
0x12b: frame_uart_px4_group_bin_0256 (RW)
0x12c: frame_uart_px4_group_bin_0032 (RW)
0x12d: frame_uart_px4_group_bin_0121 (RW)
0x12e: frame_uart_px4_group_bin_0218 (RW)
0x12f: frame_uart_px4_group_bin_0303 (RW)
0x130: frame_uart_px4_group_bin_0080 (RW)
0x131: frame_uart_px4_group_bin_0190 (RW)
0x132: frame_uart_px4_group_bin_0261 (RW)
0x134: frame_uart_px4_group_bin_0087 (RW)
0x137: frame_uart_px4_group_bin_0088 (RW)
0x13: frame_uart_px4_group_bin_0302 (RX)
0x13a: frame_uart_px4_group_bin_0233 (RW)
0x13d: frame_uart_px4_group_bin_0026 (RW)
0x140: frame_uart_px4_group_bin_0279 (RW)
0x141: frame_uart_px4_group_bin_0055 (RW)
0x142: frame_uart_px4_group_bin_0146 (RW)
0x143: frame_uart_px4_group_bin_0238 (RW)
0x146: frame_uart_px4_group_bin_0198 (RW)
0x147: frame_uart_px4_group_bin_0288 (RW)
0x148: frame_uart_px4_group_bin_0064 (RW)
0x149: frame_uart_px4_group_bin_0154 (RW)
0x14: frame_uart_px4_group_bin_0069 (RX)
0x14c: frame_uart_px4_group_bin_0111 (RW)
0x14d: frame_uart_px4_group_bin_0205 (RW)
0x14e: frame_uart_px4_group_bin_0294 (RW)
0x14f: frame_uart_px4_group_bin_0070 (RW)
0x152: frame_uart_px4_group_bin_0142 (RW)
0x153: frame_uart_px4_group_bin_0285 (RW)
0x154: frame_uart_px4_group_bin_0108 (RW)
0x155: frame_uart_px4_group_bin_0251 (RW)
0x157: frame_pilot_obj_group_bin_0009 (RWX)
0x15: frame_uart_px4_group_bin_0151 (RX)
0x16: frame_uart_px4_group_bin_0231 (RX)
0x17: frame_uart_px4_group_bin_0310 (RX)
0x18: frame_uart_px4_group_bin_0079 (RX)
0x19: frame_uart_px4_group_bin_0083 (RX)
0x1a: frame_uart_px4_group_bin_0162 (RX)
0x1b: frame_uart_px4_group_bin_0007 (RX)
0x1c: frame_uart_px4_group_bin_0089 (RX)
0x1d: frame_uart_px4_group_bin_0171 (RX)
0x1e: frame_uart_px4_group_bin_0252 (RX)
0x1f: frame_uart_px4_group_bin_0019 (RX)
0x20: frame_uart_px4_group_bin_0097 (RX)
0x30: frame_uart_px4_group_bin_0004 (RW)
0x31: frame_uart_px4_group_bin_0219 (RW)
0x32: frame_uart_px4_group_bin_0300 (RW)
0x33: frame_uart_px4_group_bin_0067 (RW)
0x34: frame_uart_px4_group_bin_0148 (RW)
0x35: frame_uart_px4_group_bin_0228 (RW)
0x36: frame_uart_px4_group_bin_0308 (RW)
0x37: frame_uart_px4_group_bin_0077 (RW)
0x38: frame_uart_px4_group_bin_0157 (RW)
0x39: frame_uart_px4_group_bin_0239 (RW)
0x3a: frame_uart_px4_group_bin_0005 (RW)
0x3b: frame_uart_px4_group_bin_0086 (RW)
0x3c: frame_uart_px4_group_bin_0169 (RW)
0x3d: frame_uart_px4_group_bin_0250 (RW)
0x3e: frame_uart_px4_group_bin_0017 (RW)
0x3f: frame_uart_px4_group_bin_0095 (RW)
0x40: frame_uart_px4_group_bin_0178 (RW)
0x41: frame_uart_px4_group_bin_0260 (RW)
0x42: frame_uart_px4_group_bin_0027 (RW)
0x43: frame_uart_px4_group_bin_0105 (RW)
0x44: frame_uart_px4_group_bin_0188 (RW)
0x45: frame_uart_px4_group_bin_0269 (RW)
0x46: frame_uart_px4_group_bin_0035 (RW)
0x47: frame_uart_px4_group_bin_0115 (RW)
0x48: frame_uart_px4_group_bin_0199 (RW)
0x49: frame_uart_px4_group_bin_0278 (RW)
0x4a: frame_uart_px4_group_bin_0044 (RW)
0x4b: frame_uart_px4_group_bin_0124 (RW)
0x4c: frame_uart_px4_group_bin_0208 (RW)
0x4d: frame_uart_px4_group_bin_0289 (RW)
0x4e: frame_uart_px4_group_bin_0054 (RW)
0x4f: frame_uart_px4_group_bin_0134 (RW)
0x50: frame_uart_px4_group_bin_0216 (RW)
0x51: frame_uart_px4_group_bin_0298 (RW)
0x52: frame_uart_px4_group_bin_0065 (RW)
0x53: frame_uart_px4_group_bin_0145 (RW)
0x54: frame_uart_px4_group_bin_0226 (RW)
0x55: frame_uart_px4_group_bin_0306 (RW)
0x56: frame_uart_px4_group_bin_0074 (RW)
0x57: frame_uart_px4_group_bin_0155 (RW)
0x58: frame_uart_px4_group_bin_0237 (RW)
0x59: frame_uart_px4_group_bin_0002 (RW)
0x5a: frame_uart_px4_group_bin_0084 (RW)
0x5b: frame_uart_px4_group_bin_0166 (RW)
0x5c: frame_uart_px4_group_bin_0247 (RW)
0x5d: frame_uart_px4_group_bin_0014 (RW)
0x5e: frame_uart_px4_group_bin_0093 (RW)
0x5f: frame_uart_px4_group_bin_0175 (RW)
0x60: frame_uart_px4_group_bin_0257 (RW)
0x61: frame_uart_px4_group_bin_0024 (RW)
0x62: frame_uart_px4_group_bin_0102 (RW)
0x63: frame_uart_px4_group_bin_0185 (RW)
0x64: frame_uart_px4_group_bin_0266 (RW)
0x65: frame_uart_px4_group_bin_0033 (RW)
0x66: frame_uart_px4_group_bin_0113 (RW)
0x67: frame_uart_px4_group_bin_0241 (RW)
0x68: frame_uart_px4_group_bin_0276 (RW)
0x69: frame_uart_px4_group_bin_0042 (RW)
0x6a: frame_uart_px4_group_bin_0122 (RW)
0x6b: frame_uart_px4_group_bin_0206 (RW)
0x6c: frame_uart_px4_group_bin_0287 (RW)
0x6d: frame_uart_px4_group_bin_0051 (RW)
0x6e: frame_uart_px4_group_bin_0131 (RW)
0x6f: frame_uart_px4_group_bin_0214 (RW)
0x70: frame_uart_px4_group_bin_0295 (RW)
0x71: frame_uart_px4_group_bin_0063 (RW)
0x72: frame_uart_px4_group_bin_0141 (RW)
0x73: frame_uart_px4_group_bin_0223 (RW)
0x74: frame_uart_px4_group_bin_0304 (RW)
0x75: frame_uart_px4_group_bin_0072 (RW)
0x76: frame_uart_px4_group_bin_0153 (RW)
0x77: frame_uart_px4_group_bin_0235 (RW)
0x78: frame_uart_px4_group_bin_0313 (RW)
0x79: frame_uart_px4_group_bin_0081 (RW)
0x7a: frame_uart_px4_group_bin_0163 (RW)
0x7b: frame_uart_px4_group_bin_0244 (RW)
0x7c: frame_uart_px4_group_bin_0011 (RW)
0x7d: frame_uart_px4_group_bin_0091 (RW)
0x7e: frame_uart_px4_group_bin_0173 (RW)
0x7f: frame_uart_px4_group_bin_0254 (RW)
0x80: frame_uart_px4_group_bin_0022 (RW)
0x81: frame_uart_px4_group_bin_0100 (RW)
0x82: frame_uart_px4_group_bin_0182 (RW)
0x83: frame_uart_px4_group_bin_0264 (RW)
0x84: frame_uart_px4_group_bin_0030 (RW)
0x85: frame_uart_px4_group_bin_0110 (RW)
0x86: frame_uart_px4_group_bin_0194 (RW)
0x87: frame_uart_px4_group_bin_0273 (RW)
0x88: frame_uart_px4_group_bin_0039 (RW)
0x89: frame_uart_px4_group_bin_0119 (RW)
0x8a: frame_uart_px4_group_bin_0204 (RW)
0x8b: frame_uart_px4_group_bin_0284 (RW)
0x8c: frame_uart_px4_group_bin_0048 (RW)
0x8d: frame_uart_px4_group_bin_0129 (RW)
0x8e: frame_uart_px4_group_bin_0212 (RW)
0x8f: frame_uart_px4_group_bin_0293 (RW)
0x90: frame_uart_px4_group_bin_0060 (RW)
0x91: frame_uart_px4_group_bin_0139 (RW)
0x92: frame_uart_px4_group_bin_0172 (RW)
0x93: frame_uart_px4_group_bin_0263 (RW)
0x94: frame_uart_px4_group_bin_0038 (RW)
0x95: frame_uart_px4_group_bin_0128 (RW)
0x96: frame_uart_px4_group_bin_0220 (RW)
0x97: frame_uart_px4_group_bin_0309 (RW)
0x98: frame_uart_px4_group_bin_0125 (RW)
0x99: frame_uart_px4_group_bin_0161 (RW)
0x9a: frame_uart_px4_group_bin_0242 (RW)
0x9b: frame_uart_px4_group_bin_0046 (RW)
0x9c: frame_uart_px4_group_bin_0136 (RW)
0x9d: frame_uart_px4_group_bin_0200 (RW)
0x9e: frame_uart_px4_group_bin_0025 (RW)
0x9f: frame_uart_px4_group_bin_0164 (RW)
0xa0: frame_uart_px4_group_bin_0189 (RW)
0xa1: frame_uart_px4_group_bin_0180 (RW)
0xa2: frame_uart_px4_group_bin_0262 (RW)
0xa3: frame_uart_px4_group_bin_0028 (RW)
0xa4: frame_uart_px4_group_bin_0107 (RW)
0xa5: frame_uart_px4_group_bin_0191 (RW)
0xa6: frame_uart_px4_group_bin_0271 (RW)
0xa7: frame_uart_px4_group_bin_0037 (RW)
0xa8: frame_uart_px4_group_bin_0117 (RW)
0xa9: frame_uart_px4_group_bin_0202 (RW)
0xaa: frame_uart_px4_group_bin_0281 (RW)
0xab: frame_uart_px4_group_bin_0246 (RW)
0xac: frame_uart_px4_group_bin_0126 (RW)
0xad: frame_uart_px4_group_bin_0210 (RW)
0xae: frame_uart_px4_group_bin_0291 (RW)
0xaf: frame_uart_px4_group_bin_0057 (RW)
0xb0: frame_uart_px4_group_bin_0071 (RW)
0xb1: frame_uart_px4_group_bin_0255 (RW)
0xb2: frame_uart_px4_group_bin_0253 (RW)
0xb3: frame_uart_px4_group_bin_0029 (RW)
0xb4: frame_uart_px4_group_bin_0118 (RW)
0xb5: frame_uart_px4_group_bin_0211 (RW)
0xb6: frame_uart_px4_group_bin_0301 (RW)
0xb7: frame_uart_px4_group_bin_0078 (RW)
0xb8: frame_uart_px4_group_bin_0217 (RW)
0xb9: frame_uart_px4_group_bin_0043 (RW)
0xba: frame_uart_px4_group_bin_0183 (RW)
0xbb: frame_uart_px4_group_bin_0008 (RW)
0xbc: frame_uart_px4_group_bin_0149 (RW)
0xbd: frame_uart_px4_group_bin_0290 (RW)
0xbe: frame_uart_px4_group_bin_0114 (RW)
0xbf: frame_uart_px4_group_bin_0009 (RW)
0xc0: frame_uart_px4_group_bin_0270 (RW)
0xc1: frame_uart_px4_group_bin_0045 (RW)
0xc2: frame_uart_px4_group_bin_0135 (RW)
0xc3: frame_uart_px4_group_bin_0227 (RW)
0xc4: frame_uart_px4_group_bin_0003 (RW)
0xc5: frame_uart_px4_group_bin_0094 (RW)
0xc6: frame_uart_px4_group_bin_0186 (RW)
0xc7: frame_uart_px4_group_bin_0277 (RW)
0xc8: frame_uart_px4_group_bin_0053 (RW)
0xc9: frame_uart_px4_group_bin_0143 (RW)
0xca: frame_uart_px4_group_bin_0236 (RW)
0xcb: frame_uart_px4_group_bin_0013 (RW)
0xcc: frame_uart_px4_group_bin_0101 (RW)
0xcd: frame_uart_px4_group_bin_0196 (RW)
0xce: frame_uart_px4_group_bin_0286 (RW)
0xcf: frame_uart_px4_group_bin_0061 (RW)
0xd0: frame_uart_px4_group_bin_0152 (RW)
0xd1: frame_uart_px4_group_bin_0243 (RW)
0xd2: frame_uart_px4_group_bin_0021 (RW)
0xd3: frame_uart_px4_group_bin_0109 (RW)
0xd4: frame_uart_px4_group_bin_0203 (RW)
0xd5: frame_uart_px4_group_bin_0292 (RW)
0xd6: frame_uart_px4_group_bin_0068 (RW)
0xd7: frame_uart_px4_group_bin_0160 (RW)
0xd8: frame_uart_px4_group_bin_0307 (RW)
0xd9: frame_uart_px4_group_bin_0132 (RW)
0xda: frame_uart_px4_group_bin_0274 (RW)
0xdb: frame_uart_px4_group_bin_0098 (RW)
0xdc: frame_uart_px4_group_bin_0240 (RW)
0xdd: frame_uart_px4_group_bin_0066 (RW)
0xde: frame_uart_px4_group_bin_0207 (RW)
0xdf: frame_uart_px4_group_bin_0031 (RW)
0xe0: frame_uart_px4_group_bin_0036 (RW)
0xe1: frame_uart_px4_group_bin_0311 (RW)
0xe2: frame_uart_px4_group_bin_0137 (RW)
0xe3: frame_uart_px4_group_bin_0280 (RW)
0xe4: frame_uart_px4_group_bin_0085 (RW)
0xe5: frame_uart_px4_group_bin_0176 (RW)
0xe6: frame_uart_px4_group_bin_0267 (RW)
0xe7: frame_uart_px4_group_bin_0197 (RW)
0xe8: frame_uart_px4_group_bin_0133 (RW)
0xe9: frame_uart_px4_group_bin_0225 (RW)
0xea: frame_uart_px4_group_bin_0096 (RW)
0xeb: frame_uart_px4_group_bin_0092 (RW)
0xec: frame_uart_px4_group_bin_0184 (RW)
0xed: frame_uart_px4_group_bin_0275 (RW)
0xee: frame_uart_px4_group_bin_0050 (RW)
0xef: frame_uart_px4_group_bin_0140 (RW)
0xf0: frame_uart_px4_group_bin_0234 (RW)
0xf1: frame_uart_px4_group_bin_0010 (RW)
0xf2: frame_uart_px4_group_bin_0099 (RW)
0xf3: frame_uart_px4_group_bin_0193 (RW)
0xf4: frame_uart_px4_group_bin_0283 (RW)
0xf5: frame_uart_px4_group_bin_0059 (RW)
0xf6: frame_uart_px4_group_bin_0150 (RW)
0xf7: frame_uart_px4_group_bin_0020 (RW)
0xf8: frame_uart_px4_group_bin_0104 (RW)
0xf9: frame_uart_px4_group_bin_0224 (RW)
0xfa: frame_uart_px4_group_bin_0049 (RW)
0xfb: frame_uart_px4_group_bin_0192 (RW)
0xfc: frame_uart_px4_group_bin_0018 (RW)
0xfd: frame_uart_px4_group_bin_0156 (RW)
0xfe: frame_uart_px4_group_bin_0296 (RW)
0xff: frame_uart_px4_group_bin_0120 (RW)
}
pt_uart_px4_group_bin_0246 {
0x0: frame_uart_px4_group_bin_0245 (RW, uncached)
}
pt_vm_group_bin_0000 {
0x100: frame_vm_group_bin_5798 (RW)
0x101: frame_vm_group_bin_22087 (RW)
0x102: frame_vm_group_bin_14936 (RW)
0x103: frame_vm_group_bin_7720 (RW)
0x104: frame_vm_group_bin_0558 (RW)
0x105: frame_vm_group_bin_16751 (RW)
0x106: frame_vm_group_bin_9542 (RW)
0x107: frame_vm_group_bin_2382 (RW)
0x108: frame_vm_group_bin_18478 (RW)
0x109: frame_vm_group_bin_11394 (RW)
0x10: frame_vm_group_bin_11624 (RX)
0x10a: frame_vm_group_bin_4209 (RW)
0x10b: frame_vm_group_bin_20305 (RW)
0x10c: frame_vm_group_bin_13110 (RW)
0x10d: frame_vm_group_bin_10444 (RW)
0x10e: frame_vm_group_bin_22118 (RW)
0x10f: frame_vm_group_bin_14969 (RW)
0x110: frame_vm_group_bin_7753 (RW)
0x111: frame_vm_group_bin_0589 (RW)
0x112: frame_vm_group_bin_16784 (RW)
0x113: frame_vm_group_bin_9575 (RW)
0x114: frame_vm_group_bin_2415 (RW)
0x115: frame_vm_group_bin_18505 (RW)
0x116: frame_vm_group_bin_11426 (RW)
0x117: frame_vm_group_bin_4242 (RW)
0x118: frame_vm_group_bin_20340 (RW)
0x119: frame_vm_group_bin_13143 (RW)
0x11: frame_vm_group_bin_22176 (RX)
0x11a: frame_vm_group_bin_15096 (RW)
0x11b: frame_vm_group_bin_22152 (RW)
0x11c: frame_vm_group_bin_15003 (RW)
0x11d: frame_vm_group_bin_7787 (RW)
0x11e: frame_vm_group_bin_9342 (RW)
0x11f: frame_vm_group_bin_16818 (RW)
0x120: frame_vm_group_bin_9609 (RW)
0x121: frame_vm_group_bin_2448 (RW)
0x122: frame_vm_group_bin_18534 (RW)
0x123: frame_vm_group_bin_11460 (RW)
0x124: frame_vm_group_bin_4276 (RW)
0x125: frame_vm_group_bin_20374 (RW)
0x126: frame_vm_group_bin_13177 (RW)
0x127: frame_vm_group_bin_19731 (RW)
0x128: frame_vm_group_bin_22185 (RW)
0x129: frame_vm_group_bin_15034 (RW)
0x12: frame_vm_group_bin_10765 (RX)
0x12a: frame_vm_group_bin_7820 (RW)
0x12b: frame_vm_group_bin_0655 (RW)
0x12c: frame_vm_group_bin_16851 (RW)
0x12d: frame_vm_group_bin_9642 (RW)
0x12e: frame_vm_group_bin_2480 (RW)
0x12f: frame_vm_group_bin_18559 (RW)
0x130: frame_vm_group_bin_11493 (RW)
0x131: frame_vm_group_bin_4309 (RW)
0x132: frame_vm_group_bin_20407 (RW)
0x133: frame_vm_group_bin_13210 (RW)
0x134: frame_vm_group_bin_1086 (RW)
0x135: frame_vm_group_bin_22218 (RW)
0x136: frame_vm_group_bin_15059 (RW)
0x137: frame_vm_group_bin_7852 (RW)
0x138: frame_vm_group_bin_0688 (RW)
0x139: frame_vm_group_bin_16883 (RW)
0x13: frame_vm_group_bin_3578 (RX)
0x13a: frame_vm_group_bin_9676 (RW)
0x13b: frame_vm_group_bin_2514 (RW)
0x13c: frame_vm_group_bin_18591 (RW)
0x13d: frame_vm_group_bin_11527 (RW)
0x13e: frame_vm_group_bin_4345 (RW)
0x13f: frame_vm_group_bin_20441 (RW)
0x140: frame_vm_group_bin_13244 (RW)
0x141: frame_vm_group_bin_6074 (RW)
0x142: frame_vm_group_bin_22252 (RW)
0x143: frame_vm_group_bin_15086 (RW)
0x144: frame_vm_group_bin_7886 (RW)
0x145: frame_vm_group_bin_0722 (RW)
0x146: frame_vm_group_bin_16916 (RW)
0x147: frame_vm_group_bin_9708 (RW)
0x148: frame_vm_group_bin_2547 (RW)
0x149: frame_vm_group_bin_18624 (RW)
0x14: frame_vm_group_bin_19680 (RX)
0x14a: frame_vm_group_bin_11558 (RW)
0x14b: frame_vm_group_bin_4378 (RW)
0x14c: frame_vm_group_bin_20474 (RW)
0x14d: frame_vm_group_bin_13277 (RW)
0x14e: frame_vm_group_bin_10469 (RW)
0x14f: frame_vm_group_bin_22284 (RW)
0x150: frame_vm_group_bin_15110 (RW)
0x151: frame_vm_group_bin_7919 (RW)
0x152: frame_vm_group_bin_0755 (RW)
0x153: frame_vm_group_bin_16949 (RW)
0x154: frame_vm_group_bin_9741 (RW)
0x155: frame_vm_group_bin_2580 (RW)
0x156: frame_vm_group_bin_18656 (RW)
0x157: frame_vm_group_bin_11585 (RW)
0x158: frame_vm_group_bin_4411 (RW)
0x159: frame_vm_group_bin_20507 (RW)
0x15: frame_vm_group_bin_12507 (RX)
0x15a: frame_vm_group_bin_13311 (RW)
0x15b: frame_vm_group_bin_6136 (RW)
0x15c: frame_vm_group_bin_22318 (RW)
0x15d: frame_vm_group_bin_15137 (RW)
0x15e: frame_vm_group_bin_7954 (RW)
0x15f: frame_vm_group_bin_0789 (RW)
0x160: frame_vm_group_bin_16983 (RW)
0x161: frame_vm_group_bin_9775 (RW)
0x162: frame_vm_group_bin_2614 (RW)
0x163: frame_vm_group_bin_18690 (RW)
0x164: frame_vm_group_bin_11613 (RW)
0x165: frame_vm_group_bin_4445 (RW)
0x166: frame_vm_group_bin_20541 (RW)
0x167: frame_vm_group_bin_13343 (RW)
0x168: frame_vm_group_bin_6168 (RW)
0x169: frame_vm_group_bin_22350 (RW)
0x16: frame_vm_group_bin_5417 (RX)
0x16a: frame_vm_group_bin_15166 (RW)
0x16b: frame_vm_group_bin_7986 (RW)
0x16c: frame_vm_group_bin_0821 (RW)
0x16d: frame_vm_group_bin_17016 (RW)
0x16e: frame_vm_group_bin_9808 (RW)
0x16f: frame_vm_group_bin_2647 (RW)
0x170: frame_vm_group_bin_18722 (RW)
0x171: frame_vm_group_bin_11635 (RW)
0x172: frame_vm_group_bin_4478 (RW)
0x173: frame_vm_group_bin_20574 (RW)
0x174: frame_vm_group_bin_13375 (RW)
0x175: frame_vm_group_bin_6199 (RW)
0x176: frame_vm_group_bin_22383 (RW)
0x177: frame_vm_group_bin_15199 (RW)
0x178: frame_vm_group_bin_8016 (RW)
0x179: frame_vm_group_bin_0854 (RW)
0x17: frame_vm_group_bin_21512 (RX)
0x17a: frame_vm_group_bin_17050 (RW)
0x17b: frame_vm_group_bin_9842 (RW)
0x17c: frame_vm_group_bin_2681 (RW)
0x17d: frame_vm_group_bin_18754 (RW)
0x17e: frame_vm_group_bin_11659 (RW)
0x17f: frame_vm_group_bin_4512 (RW)
0x180: frame_vm_group_bin_20608 (RW)
0x181: frame_vm_group_bin_13408 (RW)
0x182: frame_vm_group_bin_6227 (RW)
0x183: frame_vm_group_bin_22416 (RW)
0x184: frame_vm_group_bin_15234 (RW)
0x185: frame_vm_group_bin_8046 (RW)
0x186: frame_vm_group_bin_0888 (RW)
0x187: frame_vm_group_bin_17083 (RW)
0x188: frame_vm_group_bin_9875 (RW)
0x189: frame_vm_group_bin_2714 (RW)
0x18: frame_vm_group_bin_14336 (RX)
0x18a: frame_vm_group_bin_18787 (RW)
0x18b: frame_vm_group_bin_16234 (RW)
0x18c: frame_vm_group_bin_4545 (RW)
0x18d: frame_vm_group_bin_20641 (RW)
0x18e: frame_vm_group_bin_13441 (RW)
0x18f: frame_vm_group_bin_6257 (RW)
0x190: frame_vm_group_bin_22449 (RW)
0x191: frame_vm_group_bin_15267 (RW)
0x192: frame_vm_group_bin_8077 (RW)
0x193: frame_vm_group_bin_0921 (RW)
0x194: frame_vm_group_bin_17116 (RW)
0x195: frame_vm_group_bin_9907 (RW)
0x196: frame_vm_group_bin_2747 (RW)
0x197: frame_vm_group_bin_18820 (RW)
0x198: frame_vm_group_bin_11709 (RW)
0x199: frame_vm_group_bin_4573 (RW)
0x19: frame_vm_group_bin_7122 (RX)
0x19a: frame_vm_group_bin_20674 (RW)
0x19b: frame_vm_group_bin_13475 (RW)
0x19c: frame_vm_group_bin_6290 (RW)
0x19d: frame_vm_group_bin_22483 (RW)
0x19e: frame_vm_group_bin_15300 (RW)
0x19f: frame_vm_group_bin_8109 (RW)
0x1a0: frame_vm_group_bin_0955 (RW)
0x1a1: frame_vm_group_bin_17149 (RW)
0x1a2: frame_vm_group_bin_9939 (RW)
0x1a3: frame_vm_group_bin_2781 (RW)
0x1a4: frame_vm_group_bin_18855 (RW)
0x1a5: frame_vm_group_bin_11735 (RW)
0x1a6: frame_vm_group_bin_4598 (RW)
0x1a7: frame_vm_group_bin_20707 (RW)
0x1a8: frame_vm_group_bin_13508 (RW)
0x1a9: frame_vm_group_bin_6322 (RW)
0x1a: frame_vm_group_bin_0046 (RX)
0x1aa: frame_vm_group_bin_22516 (RW)
0x1ab: frame_vm_group_bin_15333 (RW)
0x1ac: frame_vm_group_bin_8142 (RW)
0x1ad: frame_vm_group_bin_0988 (RW)
0x1ae: frame_vm_group_bin_17181 (RW)
0x1af: frame_vm_group_bin_9972 (RW)
0x1b0: frame_vm_group_bin_2814 (RW)
0x1b1: frame_vm_group_bin_18888 (RW)
0x1b2: frame_vm_group_bin_6864 (RW)
0x1b3: frame_vm_group_bin_4622 (RW)
0x1b4: frame_vm_group_bin_20740 (RW)
0x1b5: frame_vm_group_bin_13541 (RW)
0x1b6: frame_vm_group_bin_6355 (RW)
0x1b7: frame_vm_group_bin_22548 (RW)
0x1b8: frame_vm_group_bin_15366 (RW)
0x1b9: frame_vm_group_bin_8175 (RW)
0x1b: frame_vm_group_bin_16171 (RX)
0x1ba: frame_vm_group_bin_1019 (RW)
0x1bb: frame_vm_group_bin_17213 (RW)
0x1bc: frame_vm_group_bin_10006 (RW)
0x1bd: frame_vm_group_bin_2848 (RW)
0x1be: frame_vm_group_bin_18922 (RW)
0x1bf: frame_vm_group_bin_11605 (RW)
0x1c0: frame_vm_group_bin_4653 (RW)
0x1c1: frame_vm_group_bin_20774 (RW)
0x1c2: frame_vm_group_bin_13575 (RW)
0x1c3: frame_vm_group_bin_6386 (RW)
0x1c4: frame_vm_group_bin_22582 (RW)
0x1c5: frame_vm_group_bin_15400 (RW)
0x1c6: frame_vm_group_bin_8209 (RW)
0x1c7: frame_vm_group_bin_1042 (RW)
0x1c8: frame_vm_group_bin_17245 (RW)
0x1c9: frame_vm_group_bin_10039 (RW)
0x1c: frame_vm_group_bin_8978 (RX)
0x1ca: frame_vm_group_bin_2882 (RW)
0x1cb: frame_vm_group_bin_18954 (RW)
0x1cc: frame_vm_group_bin_11811 (RW)
0x1cd: frame_vm_group_bin_4685 (RW)
0x1ce: frame_vm_group_bin_20807 (RW)
0x1cf: frame_vm_group_bin_13608 (RW)
0x1d0: frame_vm_group_bin_6418 (RW)
0x1d1: frame_vm_group_bin_22615 (RW)
0x1d2: frame_vm_group_bin_15433 (RW)
0x1d3: frame_vm_group_bin_8242 (RW)
0x1d4: frame_vm_group_bin_1063 (RW)
0x1d5: frame_vm_group_bin_17278 (RW)
0x1d6: frame_vm_group_bin_10072 (RW)
0x1d7: frame_vm_group_bin_2915 (RW)
0x1d8: frame_vm_group_bin_18985 (RW)
0x1d9: frame_vm_group_bin_20896 (RW)
0x1d: frame_vm_group_bin_1790 (RX)
0x1da: frame_vm_group_bin_4718 (RW)
0x1db: frame_vm_group_bin_20840 (RW)
0x1dc: frame_vm_group_bin_13641 (RW)
0x1dd: frame_vm_group_bin_6453 (RW)
0x1de: frame_vm_group_bin_22649 (RW)
0x1df: frame_vm_group_bin_15467 (RW)
0x1e0: frame_vm_group_bin_8275 (RW)
0x1e1: frame_vm_group_bin_1091 (RW)
0x1e2: frame_vm_group_bin_17312 (RW)
0x1e3: frame_vm_group_bin_10106 (RW)
0x1e4: frame_vm_group_bin_2949 (RW)
0x1e5: frame_vm_group_bin_19019 (RW)
0x1e6: frame_vm_group_bin_2255 (RW)
0x1e7: frame_vm_group_bin_4750 (RW)
0x1e8: frame_vm_group_bin_20865 (RW)
0x1e9: frame_vm_group_bin_13674 (RW)
0x1e: frame_vm_group_bin_17894 (RX)
0x1ea: frame_vm_group_bin_6485 (RW)
0x1eb: frame_vm_group_bin_22682 (RW)
0x1ec: frame_vm_group_bin_15500 (RW)
0x1ed: frame_vm_group_bin_8308 (RW)
0x1ee: frame_vm_group_bin_1119 (RW)
0x1ef: frame_vm_group_bin_17345 (RW)
0x1f0: frame_vm_group_bin_10139 (RW)
0x1f1: frame_vm_group_bin_2982 (RW)
0x1f2: frame_vm_group_bin_19052 (RW)
0x1f3: frame_vm_group_bin_6883 (RW)
0x1f4: frame_vm_group_bin_4783 (RW)
0x1f5: frame_vm_group_bin_20891 (RW)
0x1f6: frame_vm_group_bin_13707 (RW)
0x1f7: frame_vm_group_bin_6518 (RW)
0x1f8: frame_vm_group_bin_22715 (RW)
0x1f9: frame_vm_group_bin_15532 (RW)
0x1f: frame_vm_group_bin_10798 (RX)
0x1fa: frame_vm_group_bin_8342 (RW)
0x1fb: frame_vm_group_bin_1153 (RW)
0x1fc: frame_vm_group_bin_17378 (RW)
0x1fd: frame_vm_group_bin_10175 (RW)
0x1fe: frame_vm_group_bin_3016 (RW)
0x1ff: frame_vm_group_bin_19086 (RW)
0x20: frame_vm_group_bin_3613 (RX)
0x21: frame_vm_group_bin_19713 (RX)
0x22: frame_vm_group_bin_12541 (RX)
0x23: frame_vm_group_bin_5450 (RX)
0x24: frame_vm_group_bin_21546 (RX)
0x25: frame_vm_group_bin_14370 (RX)
0x26: frame_vm_group_bin_7155 (RX)
0x27: frame_vm_group_bin_0070 (RX)
0x28: frame_vm_group_bin_16202 (RX)
0x29: frame_vm_group_bin_9011 (RX)
0x2a: frame_vm_group_bin_1823 (RX)
0x2b: frame_vm_group_bin_17925 (RX)
0x2c: frame_vm_group_bin_10831 (RX)
0x2d: frame_vm_group_bin_3646 (RX)
0x2e: frame_vm_group_bin_19746 (RX)
0x2f: frame_vm_group_bin_12574 (RX)
0x30: frame_vm_group_bin_5482 (RX)
0x31: frame_vm_group_bin_21579 (RX)
0x32: frame_vm_group_bin_14403 (RX)
0x33: frame_vm_group_bin_7190 (RX)
0x34: frame_vm_group_bin_0097 (RX)
0x35: frame_vm_group_bin_16229 (RX)
0x36: frame_vm_group_bin_9044 (RX)
0x37: frame_vm_group_bin_1856 (RX)
0x38: frame_vm_group_bin_17956 (RX)
0x39: frame_vm_group_bin_10864 (RX)
0x3a: frame_vm_group_bin_3680 (RX)
0x3b: frame_vm_group_bin_19780 (RX)
0x3c: frame_vm_group_bin_12608 (RX)
0x3d: frame_vm_group_bin_5515 (RX)
0x3e: frame_vm_group_bin_21613 (RX)
0x3f: frame_vm_group_bin_14437 (RX)
0x40: frame_vm_group_bin_7224 (RX)
0x41: frame_vm_group_bin_0015 (RX)
0x42: frame_vm_group_bin_16258 (RX)
0x43: frame_vm_group_bin_9078 (RX)
0x44: frame_vm_group_bin_1890 (RX)
0x45: frame_vm_group_bin_17988 (RX)
0x46: frame_vm_group_bin_10898 (RX)
0x47: frame_vm_group_bin_3713 (RX)
0x48: frame_vm_group_bin_19813 (RX)
0x49: frame_vm_group_bin_12640 (RX)
0x4a: frame_vm_group_bin_5548 (RX)
0x4b: frame_vm_group_bin_21646 (RX)
0x4c: frame_vm_group_bin_14470 (RX)
0x4d: frame_vm_group_bin_7257 (RX)
0x4e: frame_vm_group_bin_4649 (RX)
0x4f: frame_vm_group_bin_16287 (RX)
0x50: frame_vm_group_bin_9111 (RX)
0x51: frame_vm_group_bin_1923 (RX)
0x52: frame_vm_group_bin_18021 (RX)
0x53: frame_vm_group_bin_10931 (RX)
0x54: frame_vm_group_bin_3746 (RX)
0x55: frame_vm_group_bin_19846 (RX)
0x65: frame_vm_group_bin_21712 (RW)
0x66: frame_vm_group_bin_14538 (RW)
0x67: frame_vm_group_bin_7323 (RW)
0x68: frame_vm_group_bin_0197 (RW)
0x69: frame_vm_group_bin_16352 (RW)
0x6a: frame_vm_group_bin_9176 (RW)
0x6b: frame_vm_group_bin_1989 (RW)
0x6c: frame_vm_group_bin_18086 (RW)
0x6d: frame_vm_group_bin_10997 (RW)
0x6e: frame_vm_group_bin_3812 (RW)
0x6f: frame_vm_group_bin_19911 (RW)
0x70: frame_vm_group_bin_12718 (RW)
0x71: frame_vm_group_bin_5645 (RW)
0x72: frame_vm_group_bin_21745 (RW)
0x73: frame_vm_group_bin_14571 (RW)
0x74: frame_vm_group_bin_7356 (RW)
0x75: frame_vm_group_bin_18565 (RW)
0x76: frame_vm_group_bin_16385 (RW)
0x77: frame_vm_group_bin_9204 (RW)
0x78: frame_vm_group_bin_2022 (RW)
0x79: frame_vm_group_bin_18118 (RW)
0x7a: frame_vm_group_bin_11031 (RW)
0x7b: frame_vm_group_bin_3846 (RW)
0x7c: frame_vm_group_bin_19944 (RW)
0x7d: frame_vm_group_bin_12744 (RW)
0x7e: frame_vm_group_bin_5679 (RW)
0x7f: frame_vm_group_bin_21778 (RW)
0x80: frame_vm_group_bin_0000 (RW)
0x81: frame_vm_group_bin_7390 (RW)
0x82: frame_vm_group_bin_0029 (RW)
0x83: frame_vm_group_bin_16419 (RW)
0x84: frame_vm_group_bin_9232 (RW)
0x85: frame_vm_group_bin_2056 (RW)
0x86: frame_vm_group_bin_18152 (RW)
0x87: frame_vm_group_bin_11064 (RW)
0x88: frame_vm_group_bin_3879 (RW)
0x89: frame_vm_group_bin_19977 (RW)
0x8a: frame_vm_group_bin_12776 (RW)
0x8b: frame_vm_group_bin_5712 (RW)
0x8c: frame_vm_group_bin_21812 (RW)
0x8d: frame_vm_group_bin_14637 (RW)
0x8e: frame_vm_group_bin_7423 (RW)
0x8f: frame_vm_group_bin_4672 (RW)
0x90: frame_vm_group_bin_16452 (RW)
0x91: frame_vm_group_bin_9255 (RW)
0x92: frame_vm_group_bin_2089 (RW)
0x93: frame_vm_group_bin_18185 (RW)
0x94: frame_vm_group_bin_11097 (RW)
0x95: frame_vm_group_bin_3912 (RW)
0x96: frame_vm_group_bin_20008 (RW)
0x97: frame_vm_group_bin_12809 (RW)
0x98: frame_vm_group_bin_5742 (RW)
0x99: frame_vm_group_bin_21845 (RW)
0x9a: frame_vm_group_bin_14671 (RW)
0x9b: frame_vm_group_bin_7457 (RW)
0x9c: frame_vm_group_bin_9298 (RW)
0x9d: frame_vm_group_bin_16486 (RW)
0x9e: frame_vm_group_bin_9281 (RW)
0x9f: frame_vm_group_bin_2124 (RW)
0xa0: frame_vm_group_bin_18218 (RW)
0xa1: frame_vm_group_bin_11130 (RW)
0xa2: frame_vm_group_bin_3945 (RW)
0xa3: frame_vm_group_bin_20042 (RW)
0xa4: frame_vm_group_bin_12842 (RW)
0xa5: frame_vm_group_bin_5768 (RW)
0xa6: frame_vm_group_bin_21879 (RW)
0xa7: frame_vm_group_bin_14704 (RW)
0xa8: frame_vm_group_bin_7490 (RW)
0xa9: frame_vm_group_bin_0336 (RW)
0xaa: frame_vm_group_bin_16519 (RW)
0xab: frame_vm_group_bin_9308 (RW)
0xac: frame_vm_group_bin_2157 (RW)
0xad: frame_vm_group_bin_18251 (RW)
0xae: frame_vm_group_bin_11163 (RW)
0xaf: frame_vm_group_bin_3978 (RW)
0xb0: frame_vm_group_bin_20075 (RW)
0xb1: frame_vm_group_bin_12875 (RW)
0xb2: frame_vm_group_bin_5791 (RW)
0xb3: frame_vm_group_bin_21912 (RW)
0xb4: frame_vm_group_bin_14736 (RW)
0xb5: frame_vm_group_bin_7522 (RW)
0xb6: frame_vm_group_bin_0368 (RW)
0xb7: frame_vm_group_bin_16552 (RW)
0xb8: frame_vm_group_bin_9340 (RW)
0xb9: frame_vm_group_bin_2189 (RW)
0xba: frame_vm_group_bin_18285 (RW)
0xbb: frame_vm_group_bin_11197 (RW)
0xbc: frame_vm_group_bin_4012 (RW)
0xbd: frame_vm_group_bin_20108 (RW)
0xbe: frame_vm_group_bin_12909 (RW)
0xbf: frame_vm_group_bin_5779 (RW)
0xc0: frame_vm_group_bin_21945 (RW)
0xc1: frame_vm_group_bin_14770 (RW)
0xc2: frame_vm_group_bin_7554 (RW)
0xc3: frame_vm_group_bin_0400 (RW)
0xc4: frame_vm_group_bin_16585 (RW)
0xc5: frame_vm_group_bin_9374 (RW)
0xc6: frame_vm_group_bin_2220 (RW)
0xc7: frame_vm_group_bin_18318 (RW)
0xc8: frame_vm_group_bin_11230 (RW)
0xc9: frame_vm_group_bin_4045 (RW)
0xca: frame_vm_group_bin_20141 (RW)
0xcb: frame_vm_group_bin_12941 (RW)
0xcc: frame_vm_group_bin_5837 (RW)
0xcd: frame_vm_group_bin_21978 (RW)
0xce: frame_vm_group_bin_14802 (RW)
0xcf: frame_vm_group_bin_7587 (RW)
0xd0: frame_vm_group_bin_0427 (RW)
0xd1: frame_vm_group_bin_16617 (RW)
0xd2: frame_vm_group_bin_9408 (RW)
0xd3: frame_vm_group_bin_2248 (RW)
0xd4: frame_vm_group_bin_18351 (RW)
0xd5: frame_vm_group_bin_11263 (RW)
0xd6: frame_vm_group_bin_4078 (RW)
0xd7: frame_vm_group_bin_20173 (RW)
0xd8: frame_vm_group_bin_12974 (RW)
0xd9: frame_vm_group_bin_5861 (RW)
0xda: frame_vm_group_bin_22011 (RW)
0xdb: frame_vm_group_bin_14836 (RW)
0xdc: frame_vm_group_bin_7621 (RW)
0xdd: frame_vm_group_bin_0461 (RW)
0xde: frame_vm_group_bin_16651 (RW)
0xdf: frame_vm_group_bin_9442 (RW)
0xe0: frame_vm_group_bin_2282 (RW)
0xe1: frame_vm_group_bin_18385 (RW)
0xe2: frame_vm_group_bin_11297 (RW)
0xe3: frame_vm_group_bin_4111 (RW)
0xe4: frame_vm_group_bin_20206 (RW)
0xe5: frame_vm_group_bin_13010 (RW)
0xe6: frame_vm_group_bin_19708 (RW)
0xe7: frame_vm_group_bin_22037 (RW)
0xe8: frame_vm_group_bin_14869 (RW)
0xe9: frame_vm_group_bin_7654 (RW)
0xea: frame_vm_group_bin_0493 (RW)
0xeb: frame_vm_group_bin_16684 (RW)
0xec: frame_vm_group_bin_9475 (RW)
0xed: frame_vm_group_bin_2315 (RW)
0xee: frame_vm_group_bin_18416 (RW)
0xef: frame_vm_group_bin_11330 (RW)
0xf0: frame_vm_group_bin_4144 (RW)
0xf1: frame_vm_group_bin_20239 (RW)
0xf2: frame_vm_group_bin_13043 (RW)
0xf3: frame_vm_group_bin_5913 (RW)
0xf4: frame_vm_group_bin_22058 (RW)
0xf5: frame_vm_group_bin_14902 (RW)
0xf6: frame_vm_group_bin_7687 (RW)
0xf7: frame_vm_group_bin_0526 (RW)
0xf8: frame_vm_group_bin_16716 (RW)
0xf9: frame_vm_group_bin_9508 (RW)
0xfa: frame_vm_group_bin_2349 (RW)
0xfb: frame_vm_group_bin_18450 (RW)
0xfc: frame_vm_group_bin_11362 (RW)
0xfd: frame_vm_group_bin_4177 (RW)
0xfe: frame_vm_group_bin_20272 (RW)
0xff: frame_vm_group_bin_13077 (RW)
}
pt_vm_group_bin_0002 {
0x0: frame_vm_group_bin_0001 (RW)
0x100: frame_vm_group_bin_7365 (RW)
0x101: frame_vm_group_bin_0235 (RW)
0x102: frame_vm_group_bin_16394 (RW)
0x103: frame_vm_group_bin_9213 (RW)
0x104: frame_vm_group_bin_2031 (RW)
0x105: frame_vm_group_bin_18127 (RW)
0x106: frame_vm_group_bin_11039 (RW)
0x107: frame_vm_group_bin_3854 (RW)
0x108: frame_vm_group_bin_19952 (RW)
0x109: frame_vm_group_bin_12751 (RW)
0x10: frame_vm_group_bin_3264 (RW)
0x10a: frame_vm_group_bin_5687 (RW)
0x10b: frame_vm_group_bin_21786 (RW)
0x10c: frame_vm_group_bin_14612 (RW)
0x10d: frame_vm_group_bin_7398 (RW)
0x10e: frame_vm_group_bin_9001 (RW)
0x10f: frame_vm_group_bin_16427 (RW)
0x110: frame_vm_group_bin_9237 (RW)
0x111: frame_vm_group_bin_2064 (RW)
0x112: frame_vm_group_bin_18160 (RW)
0x113: frame_vm_group_bin_11072 (RW)
0x114: frame_vm_group_bin_3887 (RW)
0x115: frame_vm_group_bin_19985 (RW)
0x116: frame_vm_group_bin_12784 (RW)
0x117: frame_vm_group_bin_5720 (RW)
0x118: frame_vm_group_bin_21820 (RW)
0x119: frame_vm_group_bin_14645 (RW)
0x11: frame_vm_group_bin_19334 (RW)
0x11a: frame_vm_group_bin_7432 (RW)
0x11b: frame_vm_group_bin_0282 (RW)
0x11c: frame_vm_group_bin_16461 (RW)
0x11d: frame_vm_group_bin_9261 (RW)
0x11e: frame_vm_group_bin_2098 (RW)
0x11f: frame_vm_group_bin_18193 (RW)
0x120: frame_vm_group_bin_11106 (RW)
0x121: frame_vm_group_bin_3921 (RW)
0x122: frame_vm_group_bin_20017 (RW)
0x123: frame_vm_group_bin_12817 (RW)
0x124: frame_vm_group_bin_5750 (RW)
0x125: frame_vm_group_bin_21854 (RW)
0x126: frame_vm_group_bin_14679 (RW)
0x127: frame_vm_group_bin_7465 (RW)
0x128: frame_vm_group_bin_0312 (RW)
0x129: frame_vm_group_bin_16494 (RW)
0x12: frame_vm_group_bin_20746 (RW)
0x12a: frame_vm_group_bin_9286 (RW)
0x12b: frame_vm_group_bin_2132 (RW)
0x12c: frame_vm_group_bin_18226 (RW)
0x12d: frame_vm_group_bin_11138 (RW)
0x12e: frame_vm_group_bin_3953 (RW)
0x12f: frame_vm_group_bin_20050 (RW)
0x130: frame_vm_group_bin_12850 (RW)
0x131: frame_vm_group_bin_5773 (RW)
0x132: frame_vm_group_bin_21887 (RW)
0x133: frame_vm_group_bin_14712 (RW)
0x134: frame_vm_group_bin_7498 (RW)
0x135: frame_vm_group_bin_0344 (RW)
0x136: frame_vm_group_bin_16527 (RW)
0x137: frame_vm_group_bin_9315 (RW)
0x138: frame_vm_group_bin_2165 (RW)
0x139: frame_vm_group_bin_18259 (RW)
0x13: frame_vm_group_bin_5062 (RW)
0x13a: frame_vm_group_bin_11172 (RW)
0x13b: frame_vm_group_bin_3987 (RW)
0x13c: frame_vm_group_bin_20084 (RW)
0x13d: frame_vm_group_bin_12884 (RW)
0x13e: frame_vm_group_bin_5799 (RW)
0x13f: frame_vm_group_bin_21920 (RW)
0x140: frame_vm_group_bin_14745 (RW)
0x141: frame_vm_group_bin_7530 (RW)
0x142: frame_vm_group_bin_0376 (RW)
0x143: frame_vm_group_bin_16560 (RW)
0x144: frame_vm_group_bin_9349 (RW)
0x145: frame_vm_group_bin_2198 (RW)
0x146: frame_vm_group_bin_18293 (RW)
0x147: frame_vm_group_bin_11205 (RW)
0x148: frame_vm_group_bin_4020 (RW)
0x149: frame_vm_group_bin_20116 (RW)
0x14: frame_vm_group_bin_21159 (RW)
0x14a: frame_vm_group_bin_12917 (RW)
0x14b: frame_vm_group_bin_14765 (RW)
0x14c: frame_vm_group_bin_21953 (RW)
0x14d: frame_vm_group_bin_14777 (RW)
0x14e: frame_vm_group_bin_7562 (RW)
0x14f: frame_vm_group_bin_9024 (RW)
0x150: frame_vm_group_bin_16593 (RW)
0x151: frame_vm_group_bin_9382 (RW)
0x152: frame_vm_group_bin_2227 (RW)
0x153: frame_vm_group_bin_18326 (RW)
0x154: frame_vm_group_bin_11238 (RW)
0x155: frame_vm_group_bin_4053 (RW)
0x156: frame_vm_group_bin_20149 (RW)
0x157: frame_vm_group_bin_12949 (RW)
0x158: frame_vm_group_bin_19390 (RW)
0x159: frame_vm_group_bin_21986 (RW)
0x15: frame_vm_group_bin_13982 (RW)
0x15a: frame_vm_group_bin_14811 (RW)
0x15b: frame_vm_group_bin_7596 (RW)
0x15c: frame_vm_group_bin_0436 (RW)
0x15d: frame_vm_group_bin_16626 (RW)
0x15e: frame_vm_group_bin_9417 (RW)
0x15f: frame_vm_group_bin_2257 (RW)
0x160: frame_vm_group_bin_18360 (RW)
0x161: frame_vm_group_bin_11272 (RW)
0x162: frame_vm_group_bin_4087 (RW)
0x163: frame_vm_group_bin_20181 (RW)
0x164: frame_vm_group_bin_12983 (RW)
0x165: frame_vm_group_bin_5867 (RW)
0x166: frame_vm_group_bin_22018 (RW)
0x167: frame_vm_group_bin_14844 (RW)
0x168: frame_vm_group_bin_7629 (RW)
0x169: frame_vm_group_bin_0469 (RW)
0x16: frame_vm_group_bin_6800 (RW)
0x16a: frame_vm_group_bin_16659 (RW)
0x16b: frame_vm_group_bin_9450 (RW)
0x16c: frame_vm_group_bin_2290 (RW)
0x16d: frame_vm_group_bin_18392 (RW)
0x16e: frame_vm_group_bin_11305 (RW)
0x16f: frame_vm_group_bin_4119 (RW)
0x170: frame_vm_group_bin_20214 (RW)
0x171: frame_vm_group_bin_13018 (RW)
0x172: frame_vm_group_bin_5490 (RW)
0x173: frame_vm_group_bin_22041 (RW)
0x174: frame_vm_group_bin_14877 (RW)
0x175: frame_vm_group_bin_7662 (RW)
0x176: frame_vm_group_bin_0501 (RW)
0x177: frame_vm_group_bin_16692 (RW)
0x178: frame_vm_group_bin_9483 (RW)
0x179: frame_vm_group_bin_2323 (RW)
0x17: frame_vm_group_bin_22997 (RW)
0x17a: frame_vm_group_bin_18425 (RW)
0x17b: frame_vm_group_bin_11339 (RW)
0x17c: frame_vm_group_bin_4153 (RW)
0x17d: frame_vm_group_bin_20248 (RW)
0x17e: frame_vm_group_bin_13052 (RW)
0x17f: frame_vm_group_bin_5920 (RW)
0x180: frame_vm_group_bin_22066 (RW)
0x181: frame_vm_group_bin_14911 (RW)
0x182: frame_vm_group_bin_7696 (RW)
0x183: frame_vm_group_bin_0534 (RW)
0x184: frame_vm_group_bin_16726 (RW)
0x185: frame_vm_group_bin_9517 (RW)
0x186: frame_vm_group_bin_2357 (RW)
0x187: frame_vm_group_bin_18457 (RW)
0x188: frame_vm_group_bin_11370 (RW)
0x189: frame_vm_group_bin_4185 (RW)
0x18: frame_vm_group_bin_15814 (RW)
0x18a: frame_vm_group_bin_20280 (RW)
0x18b: frame_vm_group_bin_13085 (RW)
0x18c: frame_vm_group_bin_14787 (RW)
0x18d: frame_vm_group_bin_22094 (RW)
0x18e: frame_vm_group_bin_14944 (RW)
0x18f: frame_vm_group_bin_7728 (RW)
0x190: frame_vm_group_bin_0565 (RW)
0x191: frame_vm_group_bin_16759 (RW)
0x192: frame_vm_group_bin_9550 (RW)
0x193: frame_vm_group_bin_2390 (RW)
0x194: frame_vm_group_bin_18484 (RW)
0x195: frame_vm_group_bin_11402 (RW)
0x196: frame_vm_group_bin_4217 (RW)
0x197: frame_vm_group_bin_20313 (RW)
0x198: frame_vm_group_bin_13118 (RW)
0x199: frame_vm_group_bin_5968 (RW)
0x19: frame_vm_group_bin_8621 (RW)
0x19a: frame_vm_group_bin_22127 (RW)
0x19b: frame_vm_group_bin_14978 (RW)
0x19c: frame_vm_group_bin_7762 (RW)
0x19d: frame_vm_group_bin_0598 (RW)
0x19e: frame_vm_group_bin_16793 (RW)
0x19f: frame_vm_group_bin_9584 (RW)
0x1: frame_vm_group_bin_21822 (RW)
0x1a0: frame_vm_group_bin_2423 (RW)
0x1a1: frame_vm_group_bin_18514 (RW)
0x1a2: frame_vm_group_bin_11435 (RW)
0x1a3: frame_vm_group_bin_4251 (RW)
0x1a4: frame_vm_group_bin_20349 (RW)
0x1a5: frame_vm_group_bin_13152 (RW)
0x1a6: frame_vm_group_bin_5997 (RW)
0x1a7: frame_vm_group_bin_22160 (RW)
0x1a8: frame_vm_group_bin_15011 (RW)
0x1a9: frame_vm_group_bin_7795 (RW)
0x1a: frame_vm_group_bin_1434 (RW)
0x1aa: frame_vm_group_bin_0629 (RW)
0x1ab: frame_vm_group_bin_16826 (RW)
0x1ac: frame_vm_group_bin_9617 (RW)
0x1ad: frame_vm_group_bin_2456 (RW)
0x1ae: frame_vm_group_bin_18539 (RW)
0x1af: frame_vm_group_bin_11468 (RW)
0x1b0: frame_vm_group_bin_4284 (RW)
0x1b1: frame_vm_group_bin_20382 (RW)
0x1b2: frame_vm_group_bin_13185 (RW)
0x1b3: frame_vm_group_bin_6028 (RW)
0x1b4: frame_vm_group_bin_22193 (RW)
0x1b5: frame_vm_group_bin_15039 (RW)
0x1b6: frame_vm_group_bin_7828 (RW)
0x1b7: frame_vm_group_bin_0663 (RW)
0x1b8: frame_vm_group_bin_16859 (RW)
0x1b9: frame_vm_group_bin_9650 (RW)
0x1b: frame_vm_group_bin_17585 (RW)
0x1ba: frame_vm_group_bin_2489 (RW)
0x1bb: frame_vm_group_bin_18566 (RW)
0x1bc: frame_vm_group_bin_11502 (RW)
0x1bd: frame_vm_group_bin_4318 (RW)
0x1be: frame_vm_group_bin_20416 (RW)
0x1bf: frame_vm_group_bin_13219 (RW)
0x1c0: frame_vm_group_bin_10149 (RW)
0x1c1: frame_vm_group_bin_22227 (RW)
0x1c2: frame_vm_group_bin_15067 (RW)
0x1c3: frame_vm_group_bin_7861 (RW)
0x1c4: frame_vm_group_bin_0697 (RW)
0x1c5: frame_vm_group_bin_16891 (RW)
0x1c6: frame_vm_group_bin_9683 (RW)
0x1c7: frame_vm_group_bin_2522 (RW)
0x1c8: frame_vm_group_bin_18599 (RW)
0x1c9: frame_vm_group_bin_11535 (RW)
0x1c: frame_vm_group_bin_10445 (RW)
0x1ca: frame_vm_group_bin_4353 (RW)
0x1cb: frame_vm_group_bin_20449 (RW)
0x1cc: frame_vm_group_bin_13252 (RW)
0x1cd: frame_vm_group_bin_6080 (RW)
0x1ce: frame_vm_group_bin_22260 (RW)
0x1cf: frame_vm_group_bin_15091 (RW)
0x1d0: frame_vm_group_bin_7894 (RW)
0x1d1: frame_vm_group_bin_0730 (RW)
0x1d2: frame_vm_group_bin_16924 (RW)
0x1d3: frame_vm_group_bin_9716 (RW)
0x1d4: frame_vm_group_bin_2555 (RW)
0x1d5: frame_vm_group_bin_18632 (RW)
0x1d6: frame_vm_group_bin_11565 (RW)
0x1d7: frame_vm_group_bin_4386 (RW)
0x1d8: frame_vm_group_bin_20482 (RW)
0x1d9: frame_vm_group_bin_13285 (RW)
0x1d: frame_vm_group_bin_3298 (RW)
0x1da: frame_vm_group_bin_6112 (RW)
0x1db: frame_vm_group_bin_22293 (RW)
0x1dc: frame_vm_group_bin_15119 (RW)
0x1dd: frame_vm_group_bin_7929 (RW)
0x1de: frame_vm_group_bin_0764 (RW)
0x1df: frame_vm_group_bin_16958 (RW)
0x1e0: frame_vm_group_bin_9750 (RW)
0x1e1: frame_vm_group_bin_2589 (RW)
0x1e2: frame_vm_group_bin_18665 (RW)
0x1e3: frame_vm_group_bin_11594 (RW)
0x1e4: frame_vm_group_bin_4420 (RW)
0x1e5: frame_vm_group_bin_20516 (RW)
0x1e6: frame_vm_group_bin_13318 (RW)
0x1e7: frame_vm_group_bin_6143 (RW)
0x1e8: frame_vm_group_bin_22326 (RW)
0x1e9: frame_vm_group_bin_15142 (RW)
0x1e: frame_vm_group_bin_19368 (RW)
0x1ea: frame_vm_group_bin_7962 (RW)
0x1eb: frame_vm_group_bin_0797 (RW)
0x1ec: frame_vm_group_bin_16991 (RW)
0x1ed: frame_vm_group_bin_9783 (RW)
0x1ee: frame_vm_group_bin_2622 (RW)
0x1ef: frame_vm_group_bin_18698 (RW)
0x1f0: frame_vm_group_bin_11619 (RW)
0x1f1: frame_vm_group_bin_4453 (RW)
0x1f2: frame_vm_group_bin_20549 (RW)
0x1f3: frame_vm_group_bin_13351 (RW)
0x1f4: frame_vm_group_bin_6176 (RW)
0x1f5: frame_vm_group_bin_22358 (RW)
0x1f6: frame_vm_group_bin_15174 (RW)
0x1f7: frame_vm_group_bin_7993 (RW)
0x1f8: frame_vm_group_bin_0829 (RW)
0x1f9: frame_vm_group_bin_17024 (RW)
0x1f: frame_vm_group_bin_12190 (RW)
0x1fa: frame_vm_group_bin_9817 (RW)
0x1fb: frame_vm_group_bin_2656 (RW)
0x1fc: frame_vm_group_bin_18731 (RW)
0x1fd: frame_vm_group_bin_11641 (RW)
0x1fe: frame_vm_group_bin_4487 (RW)
0x1ff: frame_vm_group_bin_20583 (RW)
0x20: frame_vm_group_bin_5097 (RW)
0x21: frame_vm_group_bin_21193 (RW)
0x22: frame_vm_group_bin_14016 (RW)
0x23: frame_vm_group_bin_6831 (RW)
0x24: frame_vm_group_bin_23030 (RW)
0x25: frame_vm_group_bin_15847 (RW)
0x26: frame_vm_group_bin_8655 (RW)
0x27: frame_vm_group_bin_1467 (RW)
0x28: frame_vm_group_bin_12466 (RW)
0x29: frame_vm_group_bin_10478 (RW)
0x2: frame_vm_group_bin_10391 (RW)
0x2a: frame_vm_group_bin_3331 (RW)
0x2b: frame_vm_group_bin_19401 (RW)
0x2c: frame_vm_group_bin_12220 (RW)
0x2d: frame_vm_group_bin_5130 (RW)
0x2e: frame_vm_group_bin_21226 (RW)
0x2f: frame_vm_group_bin_14049 (RW)
0x30: frame_vm_group_bin_6858 (RW)
0x31: frame_vm_group_bin_23063 (RW)
0x32: frame_vm_group_bin_15880 (RW)
0x33: frame_vm_group_bin_8689 (RW)
0x34: frame_vm_group_bin_1500 (RW)
0x35: frame_vm_group_bin_17640 (RW)
0x36: frame_vm_group_bin_10511 (RW)
0x37: frame_vm_group_bin_3364 (RW)
0x38: frame_vm_group_bin_19433 (RW)
0x39: frame_vm_group_bin_12252 (RW)
0x3: frame_vm_group_bin_3231 (RW)
0x3a: frame_vm_group_bin_5164 (RW)
0x3b: frame_vm_group_bin_21260 (RW)
0x3c: frame_vm_group_bin_14083 (RW)
0x3d: frame_vm_group_bin_6884 (RW)
0x3e: frame_vm_group_bin_23097 (RW)
0x3f: frame_vm_group_bin_15914 (RW)
0x40: frame_vm_group_bin_8723 (RW)
0x41: frame_vm_group_bin_1534 (RW)
0x42: frame_vm_group_bin_17674 (RW)
0x43: frame_vm_group_bin_10544 (RW)
0x44: frame_vm_group_bin_3395 (RW)
0x45: frame_vm_group_bin_19464 (RW)
0x46: frame_vm_group_bin_12286 (RW)
0x47: frame_vm_group_bin_5197 (RW)
0x48: frame_vm_group_bin_21293 (RW)
0x49: frame_vm_group_bin_14116 (RW)
0x4: frame_vm_group_bin_19301 (RW)
0x4a: frame_vm_group_bin_6907 (RW)
0x4b: frame_vm_group_bin_23130 (RW)
0x4c: frame_vm_group_bin_15947 (RW)
0x4d: frame_vm_group_bin_8756 (RW)
0x4e: frame_vm_group_bin_1567 (RW)
0x4f: frame_vm_group_bin_17702 (RW)
0x50: frame_vm_group_bin_10577 (RW)
0x51: frame_vm_group_bin_3419 (RW)
0x52: frame_vm_group_bin_19497 (RW)
0x53: frame_vm_group_bin_12319 (RW)
0x54: frame_vm_group_bin_5230 (RW)
0x55: frame_vm_group_bin_21325 (RW)
0x56: frame_vm_group_bin_14149 (RW)
0x57: frame_vm_group_bin_6937 (RW)
0x58: frame_vm_group_bin_23162 (RW)
0x59: frame_vm_group_bin_15982 (RW)
0x5: frame_vm_group_bin_12127 (RW)
0x5a: frame_vm_group_bin_8790 (RW)
0x5b: frame_vm_group_bin_1601 (RW)
0x5c: frame_vm_group_bin_17728 (RW)
0x5d: frame_vm_group_bin_10611 (RW)
0x5e: frame_vm_group_bin_3442 (RW)
0x5f: frame_vm_group_bin_19531 (RW)
0x60: frame_vm_group_bin_12352 (RW)
0x61: frame_vm_group_bin_5264 (RW)
0x62: frame_vm_group_bin_21358 (RW)
0x63: frame_vm_group_bin_14182 (RW)
0x64: frame_vm_group_bin_6969 (RW)
0x65: frame_vm_group_bin_23195 (RW)
0x66: frame_vm_group_bin_16016 (RW)
0x67: frame_vm_group_bin_8823 (RW)
0x68: frame_vm_group_bin_1634 (RW)
0x69: frame_vm_group_bin_17755 (RW)
0x6: frame_vm_group_bin_5029 (RW)
0x6a: frame_vm_group_bin_10644 (RW)
0x6b: frame_vm_group_bin_3467 (RW)
0x6c: frame_vm_group_bin_19564 (RW)
0x6d: frame_vm_group_bin_12385 (RW)
0x6e: frame_vm_group_bin_5297 (RW)
0x6f: frame_vm_group_bin_21391 (RW)
0x70: frame_vm_group_bin_14215 (RW)
0x71: frame_vm_group_bin_7002 (RW)
0x72: frame_vm_group_bin_23219 (RW)
0x73: frame_vm_group_bin_16049 (RW)
0x74: frame_vm_group_bin_8856 (RW)
0x75: frame_vm_group_bin_1667 (RW)
0x76: frame_vm_group_bin_17785 (RW)
0x77: frame_vm_group_bin_10675 (RW)
0x78: frame_vm_group_bin_3493 (RW)
0x79: frame_vm_group_bin_19598 (RW)
0x7: frame_vm_group_bin_21127 (RW)
0x7a: frame_vm_group_bin_12419 (RW)
0x7b: frame_vm_group_bin_5329 (RW)
0x7c: frame_vm_group_bin_21424 (RW)
0x7d: frame_vm_group_bin_14248 (RW)
0x7e: frame_vm_group_bin_7035 (RW)
0x7f: frame_vm_group_bin_23241 (RW)
0x80: frame_vm_group_bin_16082 (RW)
0x81: frame_vm_group_bin_8888 (RW)
0x82: frame_vm_group_bin_1700 (RW)
0x83: frame_vm_group_bin_17815 (RW)
0x84: frame_vm_group_bin_10708 (RW)
0x85: frame_vm_group_bin_3522 (RW)
0x86: frame_vm_group_bin_19631 (RW)
0x87: frame_vm_group_bin_12450 (RW)
0x88: frame_vm_group_bin_5360 (RW)
0x89: frame_vm_group_bin_21456 (RW)
0x8: frame_vm_group_bin_13949 (RW)
0x8a: frame_vm_group_bin_14280 (RW)
0x8b: frame_vm_group_bin_7066 (RW)
0x8c: frame_vm_group_bin_8952 (RW)
0x8d: frame_vm_group_bin_16114 (RW)
0x8e: frame_vm_group_bin_8920 (RW)
0x8f: frame_vm_group_bin_1732 (RW)
0x90: frame_vm_group_bin_17844 (RW)
0x91: frame_vm_group_bin_10740 (RW)
0x92: frame_vm_group_bin_3554 (RW)
0x93: frame_vm_group_bin_19659 (RW)
0x94: frame_vm_group_bin_12482 (RW)
0x95: frame_vm_group_bin_5392 (RW)
0x96: frame_vm_group_bin_21488 (RW)
0x97: frame_vm_group_bin_14311 (RW)
0x98: frame_vm_group_bin_7098 (RW)
0x99: frame_vm_group_bin_13592 (RW)
0x9: frame_vm_group_bin_6767 (RW)
0x9a: frame_vm_group_bin_16146 (RW)
0x9b: frame_vm_group_bin_8953 (RW)
0x9c: frame_vm_group_bin_1765 (RW)
0x9d: frame_vm_group_bin_17871 (RW)
0x9e: frame_vm_group_bin_10773 (RW)
0x9f: frame_vm_group_bin_3588 (RW)
0xa0: frame_vm_group_bin_19688 (RW)
0xa1: frame_vm_group_bin_12516 (RW)
0xa2: frame_vm_group_bin_5426 (RW)
0xa3: frame_vm_group_bin_21521 (RW)
0xa4: frame_vm_group_bin_14345 (RW)
0xa5: frame_vm_group_bin_7130 (RW)
0xa6: frame_vm_group_bin_18237 (RW)
0xa7: frame_vm_group_bin_16179 (RW)
0xa8: frame_vm_group_bin_8986 (RW)
0xa9: frame_vm_group_bin_1798 (RW)
0xa: frame_vm_group_bin_22964 (RW)
0xaa: frame_vm_group_bin_17901 (RW)
0xab: frame_vm_group_bin_10806 (RW)
0xac: frame_vm_group_bin_3621 (RW)
0xad: frame_vm_group_bin_19721 (RW)
0xae: frame_vm_group_bin_12549 (RW)
0xaf: frame_vm_group_bin_5458 (RW)
0xb0: frame_vm_group_bin_21554 (RW)
0xb1: frame_vm_group_bin_14378 (RW)
0xb2: frame_vm_group_bin_7163 (RW)
0xb3: frame_vm_group_bin_22977 (RW)
0xb4: frame_vm_group_bin_16209 (RW)
0xb5: frame_vm_group_bin_9019 (RW)
0xb6: frame_vm_group_bin_1831 (RW)
0xb7: frame_vm_group_bin_17933 (RW)
0xb8: frame_vm_group_bin_10839 (RW)
0xb9: frame_vm_group_bin_3654 (RW)
0xb: frame_vm_group_bin_15782 (RW)
0xba: frame_vm_group_bin_19755 (RW)
0xbb: frame_vm_group_bin_12583 (RW)
0xbc: frame_vm_group_bin_5491 (RW)
0xbd: frame_vm_group_bin_21588 (RW)
0xbe: frame_vm_group_bin_14412 (RW)
0xbf: frame_vm_group_bin_7199 (RW)
0xc0: frame_vm_group_bin_4343 (RW)
0xc1: frame_vm_group_bin_16238 (RW)
0xc2: frame_vm_group_bin_9053 (RW)
0xc3: frame_vm_group_bin_1865 (RW)
0xc4: frame_vm_group_bin_17965 (RW)
0xc5: frame_vm_group_bin_10872 (RW)
0xc6: frame_vm_group_bin_3688 (RW)
0xc7: frame_vm_group_bin_19788 (RW)
0xc8: frame_vm_group_bin_12616 (RW)
0xc9: frame_vm_group_bin_5523 (RW)
0xc: frame_vm_group_bin_8589 (RW)
0xca: frame_vm_group_bin_21621 (RW)
0xcb: frame_vm_group_bin_14445 (RW)
0xcc: frame_vm_group_bin_7232 (RW)
0xcd: frame_vm_group_bin_8977 (RW)
0xce: frame_vm_group_bin_16264 (RW)
0xcf: frame_vm_group_bin_9086 (RW)
0xd0: frame_vm_group_bin_1898 (RW)
0xd1: frame_vm_group_bin_17996 (RW)
0xd2: frame_vm_group_bin_10906 (RW)
0xd3: frame_vm_group_bin_3721 (RW)
0xd4: frame_vm_group_bin_19821 (RW)
0xd5: frame_vm_group_bin_12647 (RW)
0xd6: frame_vm_group_bin_5556 (RW)
0xd7: frame_vm_group_bin_21654 (RW)
0xd8: frame_vm_group_bin_14478 (RW)
0xd9: frame_vm_group_bin_7265 (RW)
0xd: frame_vm_group_bin_1400 (RW)
0xda: frame_vm_group_bin_13616 (RW)
0xdb: frame_vm_group_bin_16295 (RW)
0xdc: frame_vm_group_bin_9120 (RW)
0xdd: frame_vm_group_bin_1932 (RW)
0xde: frame_vm_group_bin_18030 (RW)
0xdf: frame_vm_group_bin_10940 (RW)
0xe0: frame_vm_group_bin_3755 (RW)
0xe1: frame_vm_group_bin_19855 (RW)
0xe2: frame_vm_group_bin_12675 (RW)
0xe3: frame_vm_group_bin_5589 (RW)
0xe4: frame_vm_group_bin_21687 (RW)
0xe5: frame_vm_group_bin_14513 (RW)
0xe6: frame_vm_group_bin_7298 (RW)
0xe7: frame_vm_group_bin_0173 (RW)
0xe8: frame_vm_group_bin_16327 (RW)
0xe9: frame_vm_group_bin_9152 (RW)
0xe: frame_vm_group_bin_3202 (RW)
0xea: frame_vm_group_bin_1964 (RW)
0xeb: frame_vm_group_bin_18062 (RW)
0xec: frame_vm_group_bin_10972 (RW)
0xed: frame_vm_group_bin_3787 (RW)
0xee: frame_vm_group_bin_19887 (RW)
0xef: frame_vm_group_bin_12698 (RW)
0xf0: frame_vm_group_bin_5620 (RW)
0xf1: frame_vm_group_bin_21720 (RW)
0xf2: frame_vm_group_bin_14546 (RW)
0xf3: frame_vm_group_bin_7331 (RW)
0xf4: frame_vm_group_bin_0205 (RW)
0xf5: frame_vm_group_bin_16360 (RW)
0xf6: frame_vm_group_bin_9183 (RW)
0xf7: frame_vm_group_bin_1997 (RW)
0xf8: frame_vm_group_bin_18094 (RW)
0xf9: frame_vm_group_bin_11005 (RW)
0xf: frame_vm_group_bin_10416 (RW)
0xfa: frame_vm_group_bin_3821 (RW)
0xfb: frame_vm_group_bin_19920 (RW)
0xfc: frame_vm_group_bin_12724 (RW)
0xfd: frame_vm_group_bin_5654 (RW)
0xfe: frame_vm_group_bin_21754 (RW)
0xff: frame_vm_group_bin_14580 (RW)
}
pt_vm_group_bin_0004 {
0x0: frame_vm_group_bin_8678 (RW)
0x100: frame_vm_group_bin_14700 (RW)
0x101: frame_vm_group_bin_7486 (RW)
0x102: frame_vm_group_bin_0332 (RW)
0x103: frame_vm_group_bin_16515 (RW)
0x104: frame_vm_group_bin_0064 (RW)
0x105: frame_vm_group_bin_2153 (RW)
0x106: frame_vm_group_bin_18247 (RW)
0x107: frame_vm_group_bin_11159 (RW)
0x108: frame_vm_group_bin_3974 (RW)
0x109: frame_vm_group_bin_20071 (RW)
0x10: frame_vm_group_bin_10531 (RW)
0x10a: frame_vm_group_bin_12871 (RW)
0x10b: frame_vm_group_bin_13263 (RW)
0x10c: frame_vm_group_bin_21908 (RW)
0x10d: frame_vm_group_bin_14733 (RW)
0x10e: frame_vm_group_bin_7518 (RW)
0x10f: frame_vm_group_bin_0364 (RW)
0x110: frame_vm_group_bin_16548 (RW)
0x111: frame_vm_group_bin_9336 (RW)
0x112: frame_vm_group_bin_2186 (RW)
0x113: frame_vm_group_bin_18280 (RW)
0x114: frame_vm_group_bin_11192 (RW)
0x115: frame_vm_group_bin_4007 (RW)
0x116: frame_vm_group_bin_20104 (RW)
0x117: frame_vm_group_bin_12904 (RW)
0x118: frame_vm_group_bin_5808 (RW)
0x119: frame_vm_group_bin_21940 (RW)
0x11: frame_vm_group_bin_3383 (RW)
0x11a: frame_vm_group_bin_14766 (RW)
0x11b: frame_vm_group_bin_7550 (RW)
0x11c: frame_vm_group_bin_0396 (RW)
0x11d: frame_vm_group_bin_16581 (RW)
0x11e: frame_vm_group_bin_9370 (RW)
0x11f: frame_vm_group_bin_2216 (RW)
0x120: frame_vm_group_bin_18314 (RW)
0x121: frame_vm_group_bin_11226 (RW)
0x122: frame_vm_group_bin_4041 (RW)
0x123: frame_vm_group_bin_20137 (RW)
0x124: frame_vm_group_bin_12937 (RW)
0x125: frame_vm_group_bin_5833 (RW)
0x126: frame_vm_group_bin_21974 (RW)
0x127: frame_vm_group_bin_14798 (RW)
0x128: frame_vm_group_bin_7583 (RW)
0x129: frame_vm_group_bin_0423 (RW)
0x12: frame_vm_group_bin_19452 (RW)
0x12a: frame_vm_group_bin_16613 (RW)
0x12b: frame_vm_group_bin_9404 (RW)
0x12c: frame_vm_group_bin_2244 (RW)
0x12d: frame_vm_group_bin_18347 (RW)
0x12e: frame_vm_group_bin_11259 (RW)
0x12f: frame_vm_group_bin_4074 (RW)
0x130: frame_vm_group_bin_20169 (RW)
0x131: frame_vm_group_bin_12970 (RW)
0x132: frame_vm_group_bin_5857 (RW)
0x133: frame_vm_group_bin_22007 (RW)
0x134: frame_vm_group_bin_14831 (RW)
0x135: frame_vm_group_bin_7616 (RW)
0x136: frame_vm_group_bin_0456 (RW)
0x137: frame_vm_group_bin_16646 (RW)
0x138: frame_vm_group_bin_9437 (RW)
0x139: frame_vm_group_bin_2277 (RW)
0x13: frame_vm_group_bin_12273 (RW)
0x13a: frame_vm_group_bin_18381 (RW)
0x13b: frame_vm_group_bin_11293 (RW)
0x13c: frame_vm_group_bin_12907 (RW)
0x13d: frame_vm_group_bin_20202 (RW)
0x13e: frame_vm_group_bin_13006 (RW)
0x13f: frame_vm_group_bin_5883 (RW)
0x140: frame_vm_group_bin_22035 (RW)
0x141: frame_vm_group_bin_14865 (RW)
0x142: frame_vm_group_bin_7650 (RW)
0x143: frame_vm_group_bin_0489 (RW)
0x144: frame_vm_group_bin_16680 (RW)
0x145: frame_vm_group_bin_9471 (RW)
0x146: frame_vm_group_bin_2311 (RW)
0x147: frame_vm_group_bin_18412 (RW)
0x148: frame_vm_group_bin_11326 (RW)
0x149: frame_vm_group_bin_4140 (RW)
0x14: frame_vm_group_bin_5184 (RW)
0x14a: frame_vm_group_bin_20235 (RW)
0x14b: frame_vm_group_bin_13039 (RW)
0x14c: frame_vm_group_bin_5909 (RW)
0x14d: frame_vm_group_bin_11864 (RW)
0x14e: frame_vm_group_bin_14898 (RW)
0x14f: frame_vm_group_bin_7683 (RW)
0x150: frame_vm_group_bin_0522 (RW)
0x151: frame_vm_group_bin_16712 (RW)
0x152: frame_vm_group_bin_9504 (RW)
0x153: frame_vm_group_bin_2344 (RW)
0x154: frame_vm_group_bin_18445 (RW)
0x155: frame_vm_group_bin_11357 (RW)
0x156: frame_vm_group_bin_4172 (RW)
0x157: frame_vm_group_bin_20268 (RW)
0x158: frame_vm_group_bin_13072 (RW)
0x159: frame_vm_group_bin_5934 (RW)
0x15: frame_vm_group_bin_21280 (RW)
0x15a: frame_vm_group_bin_22083 (RW)
0x15b: frame_vm_group_bin_14932 (RW)
0x15c: frame_vm_group_bin_7717 (RW)
0x15d: frame_vm_group_bin_0554 (RW)
0x15e: frame_vm_group_bin_16747 (RW)
0x15f: frame_vm_group_bin_9538 (RW)
0x160: frame_vm_group_bin_2378 (RW)
0x161: frame_vm_group_bin_18477 (RW)
0x162: frame_vm_group_bin_11390 (RW)
0x163: frame_vm_group_bin_4205 (RW)
0x164: frame_vm_group_bin_20301 (RW)
0x165: frame_vm_group_bin_13106 (RW)
0x166: frame_vm_group_bin_5957 (RW)
0x167: frame_vm_group_bin_22114 (RW)
0x168: frame_vm_group_bin_14965 (RW)
0x169: frame_vm_group_bin_7749 (RW)
0x16: frame_vm_group_bin_14103 (RW)
0x16a: frame_vm_group_bin_0585 (RW)
0x16b: frame_vm_group_bin_16780 (RW)
0x16c: frame_vm_group_bin_9571 (RW)
0x16d: frame_vm_group_bin_2411 (RW)
0x16e: frame_vm_group_bin_18502 (RW)
0x16f: frame_vm_group_bin_11422 (RW)
0x170: frame_vm_group_bin_4238 (RW)
0x171: frame_vm_group_bin_20336 (RW)
0x172: frame_vm_group_bin_13139 (RW)
0x173: frame_vm_group_bin_5986 (RW)
0x174: frame_vm_group_bin_22147 (RW)
0x175: frame_vm_group_bin_14998 (RW)
0x176: frame_vm_group_bin_7782 (RW)
0x177: frame_vm_group_bin_0618 (RW)
0x178: frame_vm_group_bin_16813 (RW)
0x179: frame_vm_group_bin_9604 (RW)
0x17: frame_vm_group_bin_13546 (RW)
0x17a: frame_vm_group_bin_2444 (RW)
0x17b: frame_vm_group_bin_18530 (RW)
0x17c: frame_vm_group_bin_11456 (RW)
0x17d: frame_vm_group_bin_4272 (RW)
0x17e: frame_vm_group_bin_20370 (RW)
0x17f: frame_vm_group_bin_13173 (RW)
0x180: frame_vm_group_bin_6017 (RW)
0x181: frame_vm_group_bin_22181 (RW)
0x182: frame_vm_group_bin_15032 (RW)
0x183: frame_vm_group_bin_7816 (RW)
0x184: frame_vm_group_bin_0651 (RW)
0x185: frame_vm_group_bin_16847 (RW)
0x186: frame_vm_group_bin_9638 (RW)
0x187: frame_vm_group_bin_2476 (RW)
0x188: frame_vm_group_bin_20508 (RW)
0x189: frame_vm_group_bin_11489 (RW)
0x18: frame_vm_group_bin_23117 (RW)
0x18a: frame_vm_group_bin_4305 (RW)
0x18b: frame_vm_group_bin_20403 (RW)
0x18c: frame_vm_group_bin_13206 (RW)
0x18d: frame_vm_group_bin_6045 (RW)
0x18e: frame_vm_group_bin_22214 (RW)
0x18f: frame_vm_group_bin_10492 (RW)
0x190: frame_vm_group_bin_7848 (RW)
0x191: frame_vm_group_bin_0684 (RW)
0x192: frame_vm_group_bin_16879 (RW)
0x193: frame_vm_group_bin_9671 (RW)
0x194: frame_vm_group_bin_2509 (RW)
0x195: frame_vm_group_bin_18586 (RW)
0x196: frame_vm_group_bin_11522 (RW)
0x197: frame_vm_group_bin_4338 (RW)
0x198: frame_vm_group_bin_20436 (RW)
0x199: frame_vm_group_bin_13239 (RW)
0x19: frame_vm_group_bin_15934 (RW)
0x19a: frame_vm_group_bin_6070 (RW)
0x19b: frame_vm_group_bin_22248 (RW)
0x19c: frame_vm_group_bin_15082 (RW)
0x19d: frame_vm_group_bin_7882 (RW)
0x19e: frame_vm_group_bin_0718 (RW)
0x19f: frame_vm_group_bin_16912 (RW)
0x1: frame_vm_group_bin_1488 (RW)
0x1a0: frame_vm_group_bin_9704 (RW)
0x1a1: frame_vm_group_bin_2543 (RW)
0x1a2: frame_vm_group_bin_18620 (RW)
0x1a3: frame_vm_group_bin_11556 (RW)
0x1a4: frame_vm_group_bin_4374 (RW)
0x1a5: frame_vm_group_bin_20470 (RW)
0x1a6: frame_vm_group_bin_13273 (RW)
0x1a7: frame_vm_group_bin_6100 (RW)
0x1a8: frame_vm_group_bin_22280 (RW)
0x1a9: frame_vm_group_bin_19779 (RW)
0x1a: frame_vm_group_bin_8744 (RW)
0x1aa: frame_vm_group_bin_7915 (RW)
0x1ab: frame_vm_group_bin_0751 (RW)
0x1ac: frame_vm_group_bin_16945 (RW)
0x1ad: frame_vm_group_bin_9737 (RW)
0x1ae: frame_vm_group_bin_2576 (RW)
0x1af: frame_vm_group_bin_18652 (RW)
0x1b0: frame_vm_group_bin_9770 (RW)
0x1b1: frame_vm_group_bin_4407 (RW)
0x1b2: frame_vm_group_bin_20503 (RW)
0x1b3: frame_vm_group_bin_13306 (RW)
0x1b4: frame_vm_group_bin_6131 (RW)
0x1b5: frame_vm_group_bin_22313 (RW)
0x1b6: frame_vm_group_bin_1127 (RW)
0x1b7: frame_vm_group_bin_7949 (RW)
0x1b8: frame_vm_group_bin_0784 (RW)
0x1b9: frame_vm_group_bin_16978 (RW)
0x1b: frame_vm_group_bin_1555 (RW)
0x1ba: frame_vm_group_bin_9771 (RW)
0x1bb: frame_vm_group_bin_2610 (RW)
0x1bc: frame_vm_group_bin_18686 (RW)
0x1bd: frame_vm_group_bin_11609 (RW)
0x1be: frame_vm_group_bin_4441 (RW)
0x1bf: frame_vm_group_bin_20537 (RW)
0x1c0: frame_vm_group_bin_13339 (RW)
0x1c1: frame_vm_group_bin_6164 (RW)
0x1c2: frame_vm_group_bin_22346 (RW)
0x1c3: frame_vm_group_bin_15162 (RW)
0x1c4: frame_vm_group_bin_7983 (RW)
0x1c5: frame_vm_group_bin_0817 (RW)
0x1c6: frame_vm_group_bin_17012 (RW)
0x1c7: frame_vm_group_bin_9804 (RW)
0x1c8: frame_vm_group_bin_2643 (RW)
0x1c9: frame_vm_group_bin_18718 (RW)
0x1c: frame_vm_group_bin_17691 (RW)
0x1ca: frame_vm_group_bin_19060 (RW)
0x1cb: frame_vm_group_bin_4474 (RW)
0x1cc: frame_vm_group_bin_20570 (RW)
0x1cd: frame_vm_group_bin_13372 (RW)
0x1ce: frame_vm_group_bin_6195 (RW)
0x1cf: frame_vm_group_bin_22379 (RW)
0x1d0: frame_vm_group_bin_15195 (RW)
0x1d1: frame_vm_group_bin_8013 (RW)
0x1d2: frame_vm_group_bin_0850 (RW)
0x1d3: frame_vm_group_bin_17045 (RW)
0x1d4: frame_vm_group_bin_9837 (RW)
0x1d5: frame_vm_group_bin_2676 (RW)
0x1d6: frame_vm_group_bin_18749 (RW)
0x1d7: frame_vm_group_bin_11654 (RW)
0x1d8: frame_vm_group_bin_4507 (RW)
0x1d9: frame_vm_group_bin_20603 (RW)
0x1d: frame_vm_group_bin_10565 (RW)
0x1da: frame_vm_group_bin_13404 (RW)
0x1db: frame_vm_group_bin_6223 (RW)
0x1dc: frame_vm_group_bin_22413 (RW)
0x1dd: frame_vm_group_bin_15230 (RW)
0x1de: frame_vm_group_bin_8042 (RW)
0x1df: frame_vm_group_bin_0884 (RW)
0x1e0: frame_vm_group_bin_17079 (RW)
0x1e1: frame_vm_group_bin_9871 (RW)
0x1e2: frame_vm_group_bin_2710 (RW)
0x1e3: frame_vm_group_bin_18783 (RW)
0x1e4: frame_vm_group_bin_11678 (RW)
0x1e5: frame_vm_group_bin_4541 (RW)
0x1e6: frame_vm_group_bin_20637 (RW)
0x1e7: frame_vm_group_bin_13437 (RW)
0x1e8: frame_vm_group_bin_6253 (RW)
0x1e9: frame_vm_group_bin_22445 (RW)
0x1e: frame_vm_group_bin_21797 (RW)
0x1ea: frame_vm_group_bin_15263 (RW)
0x1eb: frame_vm_group_bin_8073 (RW)
0x1ec: frame_vm_group_bin_0917 (RW)
0x1ed: frame_vm_group_bin_17112 (RW)
0x1ee: frame_vm_group_bin_9903 (RW)
0x1ef: frame_vm_group_bin_2743 (RW)
0x1f0: frame_vm_group_bin_18816 (RW)
0x1f1: frame_vm_group_bin_11705 (RW)
0x1f2: frame_vm_group_bin_4572 (RW)
0x1f3: frame_vm_group_bin_20669 (RW)
0x1f4: frame_vm_group_bin_13470 (RW)
0x1f5: frame_vm_group_bin_6285 (RW)
0x1f6: frame_vm_group_bin_22478 (RW)
0x1f7: frame_vm_group_bin_15295 (RW)
0x1f8: frame_vm_group_bin_8105 (RW)
0x1f9: frame_vm_group_bin_0950 (RW)
0x1f: frame_vm_group_bin_19485 (RW)
0x1fa: frame_vm_group_bin_17146 (RW)
0x1fb: frame_vm_group_bin_9936 (RW)
0x1fc: frame_vm_group_bin_2777 (RW)
0x1fd: frame_vm_group_bin_18851 (RW)
0x1fe: frame_vm_group_bin_11731 (RW)
0x1ff: frame_vm_group_bin_4595 (RW)
0x20: frame_vm_group_bin_12307 (RW)
0x21: frame_vm_group_bin_5218 (RW)
0x22: frame_vm_group_bin_21313 (RW)
0x23: frame_vm_group_bin_14137 (RW)
0x24: frame_vm_group_bin_6927 (RW)
0x25: frame_vm_group_bin_23150 (RW)
0x26: frame_vm_group_bin_15968 (RW)
0x27: frame_vm_group_bin_8777 (RW)
0x28: frame_vm_group_bin_1588 (RW)
0x29: frame_vm_group_bin_17717 (RW)
0x2: frame_vm_group_bin_17628 (RW)
0x2a: frame_vm_group_bin_10598 (RW)
0x2b: frame_vm_group_bin_8176 (RW)
0x2c: frame_vm_group_bin_19518 (RW)
0x2d: frame_vm_group_bin_12339 (RW)
0x2e: frame_vm_group_bin_5251 (RW)
0x2f: frame_vm_group_bin_21345 (RW)
0x30: frame_vm_group_bin_14170 (RW)
0x31: frame_vm_group_bin_6957 (RW)
0x32: frame_vm_group_bin_23183 (RW)
0x33: frame_vm_group_bin_16003 (RW)
0x34: frame_vm_group_bin_8810 (RW)
0x35: frame_vm_group_bin_1621 (RW)
0x36: frame_vm_group_bin_17743 (RW)
0x37: frame_vm_group_bin_10631 (RW)
0x38: frame_vm_group_bin_3457 (RW)
0x39: frame_vm_group_bin_19551 (RW)
0x3: frame_vm_group_bin_10499 (RW)
0x3a: frame_vm_group_bin_12373 (RW)
0x3b: frame_vm_group_bin_5285 (RW)
0x3c: frame_vm_group_bin_21379 (RW)
0x3d: frame_vm_group_bin_14203 (RW)
0x3e: frame_vm_group_bin_6990 (RW)
0x3f: frame_vm_group_bin_23213 (RW)
0x40: frame_vm_group_bin_16037 (RW)
0x41: frame_vm_group_bin_8844 (RW)
0x42: frame_vm_group_bin_1655 (RW)
0x43: frame_vm_group_bin_17774 (RW)
0x44: frame_vm_group_bin_10663 (RW)
0x45: frame_vm_group_bin_17535 (RW)
0x46: frame_vm_group_bin_19586 (RW)
0x47: frame_vm_group_bin_12406 (RW)
0x48: frame_vm_group_bin_5317 (RW)
0x49: frame_vm_group_bin_21412 (RW)
0x4: frame_vm_group_bin_3352 (RW)
0x4a: frame_vm_group_bin_14236 (RW)
0x4b: frame_vm_group_bin_7023 (RW)
0x4c: frame_vm_group_bin_7456 (RW)
0x4d: frame_vm_group_bin_16070 (RW)
0x4e: frame_vm_group_bin_8876 (RW)
0x4f: frame_vm_group_bin_1688 (RW)
0x50: frame_vm_group_bin_17805 (RW)
0x51: frame_vm_group_bin_10696 (RW)
0x52: frame_vm_group_bin_22199 (RW)
0x53: frame_vm_group_bin_19619 (RW)
0x54: frame_vm_group_bin_12438 (RW)
0x55: frame_vm_group_bin_5349 (RW)
0x56: frame_vm_group_bin_21444 (RW)
0x57: frame_vm_group_bin_14268 (RW)
0x58: frame_vm_group_bin_7055 (RW)
0x59: frame_vm_group_bin_0002 (RW)
0x5: frame_vm_group_bin_19421 (RW)
0x5a: frame_vm_group_bin_16103 (RW)
0x5b: frame_vm_group_bin_8909 (RW)
0x5c: frame_vm_group_bin_1721 (RW)
0x5d: frame_vm_group_bin_17834 (RW)
0x5e: frame_vm_group_bin_10729 (RW)
0x5f: frame_vm_group_bin_3543 (RW)
0x60: frame_vm_group_bin_19651 (RW)
0x61: frame_vm_group_bin_12471 (RW)
0x62: frame_vm_group_bin_5381 (RW)
0x63: frame_vm_group_bin_21477 (RW)
0x64: frame_vm_group_bin_14300 (RW)
0x65: frame_vm_group_bin_7087 (RW)
0x66: frame_vm_group_bin_16861 (RW)
0x67: frame_vm_group_bin_16134 (RW)
0x68: frame_vm_group_bin_8941 (RW)
0x69: frame_vm_group_bin_1753 (RW)
0x6: frame_vm_group_bin_12240 (RW)
0x6a: frame_vm_group_bin_17861 (RW)
0x6b: frame_vm_group_bin_10761 (RW)
0x6c: frame_vm_group_bin_3574 (RW)
0x6d: frame_vm_group_bin_6758 (RW)
0x6e: frame_vm_group_bin_12503 (RW)
0x6f: frame_vm_group_bin_5413 (RW)
0x70: frame_vm_group_bin_21508 (RW)
0x71: frame_vm_group_bin_14332 (RW)
0x72: frame_vm_group_bin_7118 (RW)
0x73: frame_vm_group_bin_0041 (RW)
0x74: frame_vm_group_bin_16166 (RW)
0x75: frame_vm_group_bin_8973 (RW)
0x76: frame_vm_group_bin_1785 (RW)
0x77: frame_vm_group_bin_17889 (RW)
0x78: frame_vm_group_bin_10793 (RW)
0x79: frame_vm_group_bin_3608 (RW)
0x7: frame_vm_group_bin_5151 (RW)
0x7a: frame_vm_group_bin_19709 (RW)
0x7b: frame_vm_group_bin_12537 (RW)
0x7c: frame_vm_group_bin_5447 (RW)
0x7d: frame_vm_group_bin_21542 (RW)
0x7e: frame_vm_group_bin_14366 (RW)
0x7f: frame_vm_group_bin_7151 (RW)
0x80: frame_vm_group_bin_0066 (RW)
0x81: frame_vm_group_bin_16200 (RW)
0x82: frame_vm_group_bin_9007 (RW)
0x83: frame_vm_group_bin_1819 (RW)
0x84: frame_vm_group_bin_17921 (RW)
0x85: frame_vm_group_bin_10827 (RW)
0x86: frame_vm_group_bin_3642 (RW)
0x87: frame_vm_group_bin_19742 (RW)
0x88: frame_vm_group_bin_12570 (RW)
0x89: frame_vm_group_bin_5478 (RW)
0x8: frame_vm_group_bin_21247 (RW)
0x8a: frame_vm_group_bin_21575 (RW)
0x8b: frame_vm_group_bin_14399 (RW)
0x8c: frame_vm_group_bin_7186 (RW)
0x8d: frame_vm_group_bin_0093 (RW)
0x8e: frame_vm_group_bin_16227 (RW)
0x8f: frame_vm_group_bin_9040 (RW)
0x90: frame_vm_group_bin_1852 (RW)
0x91: frame_vm_group_bin_17952 (RW)
0x92: frame_vm_group_bin_10860 (RW)
0x93: frame_vm_group_bin_3675 (RW)
0x94: frame_vm_group_bin_19775 (RW)
0x95: frame_vm_group_bin_12603 (RW)
0x96: frame_vm_group_bin_5511 (RW)
0x97: frame_vm_group_bin_21608 (RW)
0x98: frame_vm_group_bin_14432 (RW)
0x99: frame_vm_group_bin_7219 (RW)
0x9: frame_vm_group_bin_14070 (RW)
0x9a: frame_vm_group_bin_0119 (RW)
0x9b: frame_vm_group_bin_16254 (RW)
0x9c: frame_vm_group_bin_9074 (RW)
0x9d: frame_vm_group_bin_1886 (RW)
0x9e: frame_vm_group_bin_17984 (RW)
0x9f: frame_vm_group_bin_10894 (RW)
0xa0: frame_vm_group_bin_3709 (RW)
0xa1: frame_vm_group_bin_19809 (RW)
0xa2: frame_vm_group_bin_12637 (RW)
0xa3: frame_vm_group_bin_5544 (RW)
0xa4: frame_vm_group_bin_21642 (RW)
0xa5: frame_vm_group_bin_14466 (RW)
0xa6: frame_vm_group_bin_7253 (RW)
0xa7: frame_vm_group_bin_0140 (RW)
0xa8: frame_vm_group_bin_16283 (RW)
0xa9: frame_vm_group_bin_9107 (RW)
0xa: frame_vm_group_bin_8907 (RW)
0xaa: frame_vm_group_bin_1919 (RW)
0xab: frame_vm_group_bin_18017 (RW)
0xac: frame_vm_group_bin_10927 (RW)
0xad: frame_vm_group_bin_3742 (RW)
0xae: frame_vm_group_bin_19842 (RW)
0xaf: frame_vm_group_bin_12666 (RW)
0xb0: frame_vm_group_bin_5577 (RW)
0xb1: frame_vm_group_bin_21675 (RW)
0xb2: frame_vm_group_bin_14499 (RW)
0xb3: frame_vm_group_bin_7286 (RW)
0xb4: frame_vm_group_bin_0162 (RW)
0xb5: frame_vm_group_bin_16315 (RW)
0xb6: frame_vm_group_bin_9140 (RW)
0xb7: frame_vm_group_bin_1952 (RW)
0xb8: frame_vm_group_bin_18050 (RW)
0xb9: frame_vm_group_bin_10960 (RW)
0xb: frame_vm_group_bin_23084 (RW)
0xba: frame_vm_group_bin_3776 (RW)
0xbb: frame_vm_group_bin_19876 (RW)
0xbc: frame_vm_group_bin_12690 (RW)
0xbd: frame_vm_group_bin_5610 (RW)
0xbe: frame_vm_group_bin_21708 (RW)
0xbf: frame_vm_group_bin_14534 (RW)
0xc0: frame_vm_group_bin_7319 (RW)
0xc1: frame_vm_group_bin_0193 (RW)
0xc2: frame_vm_group_bin_16348 (RW)
0xc3: frame_vm_group_bin_9172 (RW)
0xc4: frame_vm_group_bin_1985 (RW)
0xc5: frame_vm_group_bin_18082 (RW)
0xc6: frame_vm_group_bin_10993 (RW)
0xc7: frame_vm_group_bin_3808 (RW)
0xc8: frame_vm_group_bin_19907 (RW)
0xc9: frame_vm_group_bin_14719 (RW)
0xc: frame_vm_group_bin_15901 (RW)
0xca: frame_vm_group_bin_5641 (RW)
0xcb: frame_vm_group_bin_21741 (RW)
0xcc: frame_vm_group_bin_14567 (RW)
0xcd: frame_vm_group_bin_7352 (RW)
0xce: frame_vm_group_bin_0224 (RW)
0xcf: frame_vm_group_bin_16381 (RW)
0xd0: frame_vm_group_bin_9203 (RW)
0xd1: frame_vm_group_bin_2018 (RW)
0xd2: frame_vm_group_bin_18114 (RW)
0xd3: frame_vm_group_bin_11026 (RW)
0xd4: frame_vm_group_bin_3841 (RW)
0xd5: frame_vm_group_bin_19939 (RW)
0xd6: frame_vm_group_bin_19342 (RW)
0xd7: frame_vm_group_bin_5674 (RW)
0xd8: frame_vm_group_bin_21774 (RW)
0xd9: frame_vm_group_bin_14600 (RW)
0xd: frame_vm_group_bin_8710 (RW)
0xda: frame_vm_group_bin_7386 (RW)
0xdb: frame_vm_group_bin_0248 (RW)
0xdc: frame_vm_group_bin_16415 (RW)
0xdd: frame_vm_group_bin_9228 (RW)
0xde: frame_vm_group_bin_2052 (RW)
0xdf: frame_vm_group_bin_18148 (RW)
0xe0: frame_vm_group_bin_11060 (RW)
0xe1: frame_vm_group_bin_3875 (RW)
0xe2: frame_vm_group_bin_19973 (RW)
0xe3: frame_vm_group_bin_12772 (RW)
0xe4: frame_vm_group_bin_5708 (RW)
0xe5: frame_vm_group_bin_21808 (RW)
0xe6: frame_vm_group_bin_14633 (RW)
0xe7: frame_vm_group_bin_7419 (RW)
0xe8: frame_vm_group_bin_0271 (RW)
0xe9: frame_vm_group_bin_16448 (RW)
0xe: frame_vm_group_bin_1521 (RW)
0xea: frame_vm_group_bin_13987 (RW)
0xeb: frame_vm_group_bin_2085 (RW)
0xec: frame_vm_group_bin_18181 (RW)
0xed: frame_vm_group_bin_11093 (RW)
0xee: frame_vm_group_bin_3908 (RW)
0xef: frame_vm_group_bin_20004 (RW)
0xf0: frame_vm_group_bin_12805 (RW)
0xf1: frame_vm_group_bin_5740 (RW)
0xf2: frame_vm_group_bin_21841 (RW)
0xf3: frame_vm_group_bin_14666 (RW)
0xf4: frame_vm_group_bin_7452 (RW)
0xf5: frame_vm_group_bin_0300 (RW)
0xf6: frame_vm_group_bin_16481 (RW)
0xf7: frame_vm_group_bin_9276 (RW)
0xf8: frame_vm_group_bin_2118 (RW)
0xf9: frame_vm_group_bin_18213 (RW)
0xf: frame_vm_group_bin_17661 (RW)
0xfa: frame_vm_group_bin_11126 (RW)
0xfb: frame_vm_group_bin_3941 (RW)
0xfc: frame_vm_group_bin_20038 (RW)
0xfd: frame_vm_group_bin_12838 (RW)
0xfe: frame_vm_group_bin_8622 (RW)
0xff: frame_vm_group_bin_21875 (RW)
}
pt_vm_group_bin_0006 {
0x0: frame_vm_group_bin_0003 (RW)
0x100: frame_vm_group_bin_11764 (RW)
0x101: frame_vm_group_bin_4366 (RW)
0x102: frame_vm_group_bin_20751 (RW)
0x103: frame_vm_group_bin_13552 (RW)
0x104: frame_vm_group_bin_6366 (RW)
0x105: frame_vm_group_bin_22559 (RW)
0x106: frame_vm_group_bin_15377 (RW)
0x107: frame_vm_group_bin_8186 (RW)
0x108: frame_vm_group_bin_1027 (RW)
0x109: frame_vm_group_bin_17223 (RW)
0x10: frame_vm_group_bin_7564 (RW)
0x10a: frame_vm_group_bin_10016 (RW)
0x10b: frame_vm_group_bin_2857 (RW)
0x10c: frame_vm_group_bin_18932 (RW)
0x10d: frame_vm_group_bin_11789 (RW)
0x10e: frame_vm_group_bin_4663 (RW)
0x10f: frame_vm_group_bin_20784 (RW)
0x110: frame_vm_group_bin_13585 (RW)
0x111: frame_vm_group_bin_6396 (RW)
0x112: frame_vm_group_bin_22592 (RW)
0x113: frame_vm_group_bin_15410 (RW)
0x114: frame_vm_group_bin_8219 (RW)
0x115: frame_vm_group_bin_22269 (RW)
0x116: frame_vm_group_bin_17255 (RW)
0x117: frame_vm_group_bin_10049 (RW)
0x118: frame_vm_group_bin_2892 (RW)
0x119: frame_vm_group_bin_16554 (RW)
0x11: frame_vm_group_bin_0406 (RW)
0x11a: frame_vm_group_bin_11822 (RW)
0x11b: frame_vm_group_bin_4696 (RW)
0x11c: frame_vm_group_bin_20818 (RW)
0x11d: frame_vm_group_bin_13619 (RW)
0x11e: frame_vm_group_bin_6429 (RW)
0x11f: frame_vm_group_bin_22626 (RW)
0x120: frame_vm_group_bin_15444 (RW)
0x121: frame_vm_group_bin_8253 (RW)
0x122: frame_vm_group_bin_3632 (RW)
0x123: frame_vm_group_bin_17289 (RW)
0x124: frame_vm_group_bin_10083 (RW)
0x125: frame_vm_group_bin_2926 (RW)
0x126: frame_vm_group_bin_18996 (RW)
0x127: frame_vm_group_bin_11852 (RW)
0x128: frame_vm_group_bin_4727 (RW)
0x129: frame_vm_group_bin_20848 (RW)
0x12: frame_vm_group_bin_16595 (RW)
0x12a: frame_vm_group_bin_13651 (RW)
0x12b: frame_vm_group_bin_6462 (RW)
0x12c: frame_vm_group_bin_22659 (RW)
0x12d: frame_vm_group_bin_15477 (RW)
0x12e: frame_vm_group_bin_8285 (RW)
0x12f: frame_vm_group_bin_8271 (RW)
0x130: frame_vm_group_bin_17322 (RW)
0x131: frame_vm_group_bin_10116 (RW)
0x132: frame_vm_group_bin_2959 (RW)
0x133: frame_vm_group_bin_19029 (RW)
0x134: frame_vm_group_bin_11880 (RW)
0x135: frame_vm_group_bin_4760 (RW)
0x136: frame_vm_group_bin_20872 (RW)
0x137: frame_vm_group_bin_13684 (RW)
0x138: frame_vm_group_bin_6495 (RW)
0x139: frame_vm_group_bin_22692 (RW)
0x13: frame_vm_group_bin_9384 (RW)
0x13a: frame_vm_group_bin_15511 (RW)
0x13b: frame_vm_group_bin_8319 (RW)
0x13c: frame_vm_group_bin_1130 (RW)
0x13d: frame_vm_group_bin_17356 (RW)
0x13e: frame_vm_group_bin_10152 (RW)
0x13f: frame_vm_group_bin_2993 (RW)
0x140: frame_vm_group_bin_19063 (RW)
0x141: frame_vm_group_bin_11904 (RW)
0x142: frame_vm_group_bin_4794 (RW)
0x143: frame_vm_group_bin_2941 (RW)
0x144: frame_vm_group_bin_13717 (RW)
0x145: frame_vm_group_bin_6529 (RW)
0x146: frame_vm_group_bin_22726 (RW)
0x147: frame_vm_group_bin_15542 (RW)
0x148: frame_vm_group_bin_8352 (RW)
0x149: frame_vm_group_bin_1163 (RW)
0x14: frame_vm_group_bin_17831 (RW)
0x14a: frame_vm_group_bin_17387 (RW)
0x14b: frame_vm_group_bin_10185 (RW)
0x14c: frame_vm_group_bin_3026 (RW)
0x14d: frame_vm_group_bin_19096 (RW)
0x14e: frame_vm_group_bin_11934 (RW)
0x14f: frame_vm_group_bin_4826 (RW)
0x150: frame_vm_group_bin_20927 (RW)
0x151: frame_vm_group_bin_13750 (RW)
0x152: frame_vm_group_bin_6562 (RW)
0x153: frame_vm_group_bin_22758 (RW)
0x154: frame_vm_group_bin_15575 (RW)
0x155: frame_vm_group_bin_8385 (RW)
0x156: frame_vm_group_bin_1196 (RW)
0x157: frame_vm_group_bin_17413 (RW)
0x158: frame_vm_group_bin_10218 (RW)
0x159: frame_vm_group_bin_3059 (RW)
0x15: frame_vm_group_bin_18328 (RW)
0x15a: frame_vm_group_bin_19129 (RW)
0x15b: frame_vm_group_bin_11965 (RW)
0x15c: frame_vm_group_bin_4860 (RW)
0x15d: frame_vm_group_bin_20955 (RW)
0x15e: frame_vm_group_bin_13785 (RW)
0x15f: frame_vm_group_bin_6596 (RW)
0x160: frame_vm_group_bin_22792 (RW)
0x161: frame_vm_group_bin_15609 (RW)
0x162: frame_vm_group_bin_8419 (RW)
0x163: frame_vm_group_bin_1230 (RW)
0x164: frame_vm_group_bin_2211 (RW)
0x165: frame_vm_group_bin_10252 (RW)
0x166: frame_vm_group_bin_3093 (RW)
0x167: frame_vm_group_bin_19161 (RW)
0x168: frame_vm_group_bin_11997 (RW)
0x169: frame_vm_group_bin_4893 (RW)
0x16: frame_vm_group_bin_11240 (RW)
0x16a: frame_vm_group_bin_20986 (RW)
0x16b: frame_vm_group_bin_13817 (RW)
0x16c: frame_vm_group_bin_6629 (RW)
0x16d: frame_vm_group_bin_22825 (RW)
0x16e: frame_vm_group_bin_15642 (RW)
0x16f: frame_vm_group_bin_8452 (RW)
0x170: frame_vm_group_bin_1262 (RW)
0x171: frame_vm_group_bin_12277 (RW)
0x172: frame_vm_group_bin_10285 (RW)
0x173: frame_vm_group_bin_3125 (RW)
0x174: frame_vm_group_bin_19194 (RW)
0x175: frame_vm_group_bin_12028 (RW)
0x176: frame_vm_group_bin_4925 (RW)
0x177: frame_vm_group_bin_21019 (RW)
0x178: frame_vm_group_bin_13846 (RW)
0x179: frame_vm_group_bin_6662 (RW)
0x17: frame_vm_group_bin_4055 (RW)
0x17a: frame_vm_group_bin_22859 (RW)
0x17b: frame_vm_group_bin_15676 (RW)
0x17c: frame_vm_group_bin_8486 (RW)
0x17d: frame_vm_group_bin_1294 (RW)
0x17e: frame_vm_group_bin_11588 (RW)
0x17f: frame_vm_group_bin_10319 (RW)
0x180: frame_vm_group_bin_3159 (RW)
0x181: frame_vm_group_bin_19228 (RW)
0x182: frame_vm_group_bin_12056 (RW)
0x183: frame_vm_group_bin_4957 (RW)
0x184: frame_vm_group_bin_21054 (RW)
0x185: frame_vm_group_bin_1483 (RW)
0x186: frame_vm_group_bin_6696 (RW)
0x187: frame_vm_group_bin_22892 (RW)
0x188: frame_vm_group_bin_15709 (RW)
0x189: frame_vm_group_bin_8518 (RW)
0x18: frame_vm_group_bin_20151 (RW)
0x18a: frame_vm_group_bin_1326 (RW)
0x18b: frame_vm_group_bin_17505 (RW)
0x18c: frame_vm_group_bin_10352 (RW)
0x18d: frame_vm_group_bin_3192 (RW)
0x18e: frame_vm_group_bin_19261 (RW)
0x18f: frame_vm_group_bin_12088 (RW)
0x190: frame_vm_group_bin_4989 (RW)
0x191: frame_vm_group_bin_21087 (RW)
0x192: frame_vm_group_bin_13909 (RW)
0x193: frame_vm_group_bin_6728 (RW)
0x194: frame_vm_group_bin_22925 (RW)
0x195: frame_vm_group_bin_15742 (RW)
0x196: frame_vm_group_bin_8550 (RW)
0x197: frame_vm_group_bin_1359 (RW)
0x198: frame_vm_group_bin_17533 (RW)
0x199: frame_vm_group_bin_10384 (RW)
0x19: frame_vm_group_bin_12951 (RW)
0x19a: frame_vm_group_bin_3226 (RW)
0x19b: frame_vm_group_bin_19295 (RW)
0x19c: frame_vm_group_bin_12121 (RW)
0x19d: frame_vm_group_bin_5023 (RW)
0x19e: frame_vm_group_bin_21121 (RW)
0x19f: frame_vm_group_bin_13943 (RW)
0x1: frame_vm_group_bin_21922 (RW)
0x1a0: frame_vm_group_bin_6761 (RW)
0x1a1: frame_vm_group_bin_22958 (RW)
0x1a2: frame_vm_group_bin_15776 (RW)
0x1a3: frame_vm_group_bin_8583 (RW)
0x1a4: frame_vm_group_bin_1394 (RW)
0x1a5: frame_vm_group_bin_2233 (RW)
0x1a6: frame_vm_group_bin_0786 (RW)
0x1a7: frame_vm_group_bin_3258 (RW)
0x1a8: frame_vm_group_bin_19328 (RW)
0x1a9: frame_vm_group_bin_12154 (RW)
0x1a: frame_vm_group_bin_9260 (RW)
0x1aa: frame_vm_group_bin_5056 (RW)
0x1ab: frame_vm_group_bin_21153 (RW)
0x1ac: frame_vm_group_bin_13976 (RW)
0x1ad: frame_vm_group_bin_6794 (RW)
0x1ae: frame_vm_group_bin_22991 (RW)
0x1af: frame_vm_group_bin_15808 (RW)
0x1b0: frame_vm_group_bin_8615 (RW)
0x1b1: frame_vm_group_bin_1427 (RW)
0x1b2: frame_vm_group_bin_17578 (RW)
0x1b3: frame_vm_group_bin_5514 (RW)
0x1b4: frame_vm_group_bin_3291 (RW)
0x1b5: frame_vm_group_bin_19361 (RW)
0x1b6: frame_vm_group_bin_12184 (RW)
0x1b7: frame_vm_group_bin_5090 (RW)
0x1b8: frame_vm_group_bin_21186 (RW)
0x1b9: frame_vm_group_bin_14009 (RW)
0x1b: frame_vm_group_bin_21989 (RW)
0x1ba: frame_vm_group_bin_6825 (RW)
0x1bb: frame_vm_group_bin_23024 (RW)
0x1bc: frame_vm_group_bin_15841 (RW)
0x1bd: frame_vm_group_bin_8649 (RW)
0x1be: frame_vm_group_bin_1461 (RW)
0x1bf: frame_vm_group_bin_17603 (RW)
0x1c0: frame_vm_group_bin_10472 (RW)
0x1c1: frame_vm_group_bin_3325 (RW)
0x1c2: frame_vm_group_bin_19395 (RW)
0x1c3: frame_vm_group_bin_12214 (RW)
0x1c4: frame_vm_group_bin_5124 (RW)
0x1c5: frame_vm_group_bin_21220 (RW)
0x1c6: frame_vm_group_bin_14043 (RW)
0x1c7: frame_vm_group_bin_6854 (RW)
0x1c8: frame_vm_group_bin_23057 (RW)
0x1c9: frame_vm_group_bin_15874 (RW)
0x1c: frame_vm_group_bin_14813 (RW)
0x1ca: frame_vm_group_bin_8683 (RW)
0x1cb: frame_vm_group_bin_1494 (RW)
0x1cc: frame_vm_group_bin_17634 (RW)
0x1cd: frame_vm_group_bin_10505 (RW)
0x1ce: frame_vm_group_bin_3358 (RW)
0x1cf: frame_vm_group_bin_19427 (RW)
0x1d0: frame_vm_group_bin_12246 (RW)
0x1d1: frame_vm_group_bin_5157 (RW)
0x1d2: frame_vm_group_bin_21253 (RW)
0x1d3: frame_vm_group_bin_14076 (RW)
0x1d4: frame_vm_group_bin_4789 (RW)
0x1d5: frame_vm_group_bin_23090 (RW)
0x1d6: frame_vm_group_bin_15907 (RW)
0x1d7: frame_vm_group_bin_8716 (RW)
0x1d8: frame_vm_group_bin_1527 (RW)
0x1d9: frame_vm_group_bin_17667 (RW)
0x1d: frame_vm_group_bin_7598 (RW)
0x1da: frame_vm_group_bin_10538 (RW)
0x1db: frame_vm_group_bin_3389 (RW)
0x1dc: frame_vm_group_bin_19458 (RW)
0x1dd: frame_vm_group_bin_12280 (RW)
0x1de: frame_vm_group_bin_5191 (RW)
0x1df: frame_vm_group_bin_21287 (RW)
0x1e0: frame_vm_group_bin_14110 (RW)
0x1e1: frame_vm_group_bin_9416 (RW)
0x1e2: frame_vm_group_bin_23124 (RW)
0x1e3: frame_vm_group_bin_15941 (RW)
0x1e4: frame_vm_group_bin_8750 (RW)
0x1e5: frame_vm_group_bin_1561 (RW)
0x1e6: frame_vm_group_bin_17696 (RW)
0x1e7: frame_vm_group_bin_10571 (RW)
0x1e8: frame_vm_group_bin_3416 (RW)
0x1e9: frame_vm_group_bin_19491 (RW)
0x1e: frame_vm_group_bin_0438 (RW)
0x1ea: frame_vm_group_bin_12313 (RW)
0x1eb: frame_vm_group_bin_5224 (RW)
0x1ec: frame_vm_group_bin_21319 (RW)
0x1ed: frame_vm_group_bin_14143 (RW)
0x1ee: frame_vm_group_bin_14082 (RW)
0x1ef: frame_vm_group_bin_23156 (RW)
0x1f0: frame_vm_group_bin_15974 (RW)
0x1f1: frame_vm_group_bin_8783 (RW)
0x1f2: frame_vm_group_bin_1594 (RW)
0x1f3: frame_vm_group_bin_17721 (RW)
0x1f4: frame_vm_group_bin_10604 (RW)
0x1f5: frame_vm_group_bin_4082 (RW)
0x1f6: frame_vm_group_bin_19524 (RW)
0x1f7: frame_vm_group_bin_12345 (RW)
0x1f8: frame_vm_group_bin_5257 (RW)
0x1f9: frame_vm_group_bin_21351 (RW)
0x1f: frame_vm_group_bin_16628 (RW)
0x1fa: frame_vm_group_bin_14177 (RW)
0x1fb: frame_vm_group_bin_6964 (RW)
0x1fc: frame_vm_group_bin_23189 (RW)
0x1fd: frame_vm_group_bin_16010 (RW)
0x1fe: frame_vm_group_bin_8817 (RW)
0x1ff: frame_vm_group_bin_1628 (RW)
0x20: frame_vm_group_bin_9419 (RW)
0x21: frame_vm_group_bin_2259 (RW)
0x22: frame_vm_group_bin_18362 (RW)
0x23: frame_vm_group_bin_11274 (RW)
0x24: frame_vm_group_bin_4089 (RW)
0x25: frame_vm_group_bin_20183 (RW)
0x26: frame_vm_group_bin_12985 (RW)
0x27: frame_vm_group_bin_5868 (RW)
0x28: frame_vm_group_bin_22020 (RW)
0x29: frame_vm_group_bin_14846 (RW)
0x2: frame_vm_group_bin_14747 (RW)
0x2a: frame_vm_group_bin_7631 (RW)
0x2b: frame_vm_group_bin_0471 (RW)
0x2c: frame_vm_group_bin_16661 (RW)
0x2d: frame_vm_group_bin_9452 (RW)
0x2e: frame_vm_group_bin_2292 (RW)
0x2f: frame_vm_group_bin_18394 (RW)
0x30: frame_vm_group_bin_11307 (RW)
0x31: frame_vm_group_bin_4121 (RW)
0x32: frame_vm_group_bin_20216 (RW)
0x33: frame_vm_group_bin_13020 (RW)
0x34: frame_vm_group_bin_18545 (RW)
0x35: frame_vm_group_bin_22043 (RW)
0x36: frame_vm_group_bin_14879 (RW)
0x37: frame_vm_group_bin_7664 (RW)
0x38: frame_vm_group_bin_0503 (RW)
0x39: frame_vm_group_bin_16694 (RW)
0x3: frame_vm_group_bin_7532 (RW)
0x3a: frame_vm_group_bin_9486 (RW)
0x3b: frame_vm_group_bin_2326 (RW)
0x3c: frame_vm_group_bin_18427 (RW)
0x3d: frame_vm_group_bin_11341 (RW)
0x3e: frame_vm_group_bin_4155 (RW)
0x3f: frame_vm_group_bin_20250 (RW)
0x40: frame_vm_group_bin_13054 (RW)
0x41: frame_vm_group_bin_5921 (RW)
0x42: frame_vm_group_bin_21846 (RW)
0x43: frame_vm_group_bin_14913 (RW)
0x44: frame_vm_group_bin_7698 (RW)
0x45: frame_vm_group_bin_0536 (RW)
0x46: frame_vm_group_bin_16728 (RW)
0x47: frame_vm_group_bin_9519 (RW)
0x48: frame_vm_group_bin_2359 (RW)
0x49: frame_vm_group_bin_18459 (RW)
0x4: frame_vm_group_bin_0378 (RW)
0x4a: frame_vm_group_bin_11372 (RW)
0x4b: frame_vm_group_bin_4187 (RW)
0x4c: frame_vm_group_bin_20282 (RW)
0x4d: frame_vm_group_bin_13087 (RW)
0x4e: frame_vm_group_bin_5943 (RW)
0x4f: frame_vm_group_bin_3225 (RW)
0x50: frame_vm_group_bin_14946 (RW)
0x51: frame_vm_group_bin_7730 (RW)
0x52: frame_vm_group_bin_0567 (RW)
0x53: frame_vm_group_bin_16761 (RW)
0x54: frame_vm_group_bin_9552 (RW)
0x55: frame_vm_group_bin_2392 (RW)
0x56: frame_vm_group_bin_18486 (RW)
0x57: frame_vm_group_bin_11404 (RW)
0x58: frame_vm_group_bin_4219 (RW)
0x59: frame_vm_group_bin_20317 (RW)
0x5: frame_vm_group_bin_16562 (RW)
0x5a: frame_vm_group_bin_13121 (RW)
0x5b: frame_vm_group_bin_9279 (RW)
0x5c: frame_vm_group_bin_22129 (RW)
0x5d: frame_vm_group_bin_14980 (RW)
0x5e: frame_vm_group_bin_7764 (RW)
0x5f: frame_vm_group_bin_0600 (RW)
0x60: frame_vm_group_bin_16795 (RW)
0x61: frame_vm_group_bin_9586 (RW)
0x62: frame_vm_group_bin_2425 (RW)
0x63: frame_vm_group_bin_18516 (RW)
0x64: frame_vm_group_bin_11437 (RW)
0x65: frame_vm_group_bin_4253 (RW)
0x66: frame_vm_group_bin_20351 (RW)
0x67: frame_vm_group_bin_13154 (RW)
0x68: frame_vm_group_bin_5999 (RW)
0x69: frame_vm_group_bin_22162 (RW)
0x6: frame_vm_group_bin_9351 (RW)
0x6a: frame_vm_group_bin_15013 (RW)
0x6b: frame_vm_group_bin_7797 (RW)
0x6c: frame_vm_group_bin_0631 (RW)
0x6d: frame_vm_group_bin_16828 (RW)
0x6e: frame_vm_group_bin_9619 (RW)
0x6f: frame_vm_group_bin_2458 (RW)
0x70: frame_vm_group_bin_2488 (RW)
0x71: frame_vm_group_bin_11470 (RW)
0x72: frame_vm_group_bin_4286 (RW)
0x73: frame_vm_group_bin_20384 (RW)
0x74: frame_vm_group_bin_13187 (RW)
0x75: frame_vm_group_bin_6030 (RW)
0x76: frame_vm_group_bin_22195 (RW)
0x77: frame_vm_group_bin_15041 (RW)
0x78: frame_vm_group_bin_7830 (RW)
0x79: frame_vm_group_bin_0665 (RW)
0x7: frame_vm_group_bin_2200 (RW)
0x7a: frame_vm_group_bin_16862 (RW)
0x7b: frame_vm_group_bin_9653 (RW)
0x7c: frame_vm_group_bin_2491 (RW)
0x7d: frame_vm_group_bin_18568 (RW)
0x7e: frame_vm_group_bin_11504 (RW)
0x7f: frame_vm_group_bin_4320 (RW)
0x80: frame_vm_group_bin_20418 (RW)
0x81: frame_vm_group_bin_13221 (RW)
0x82: frame_vm_group_bin_6056 (RW)
0x83: frame_vm_group_bin_22229 (RW)
0x84: frame_vm_group_bin_20415 (RW)
0x85: frame_vm_group_bin_7863 (RW)
0x86: frame_vm_group_bin_0699 (RW)
0x87: frame_vm_group_bin_16893 (RW)
0x88: frame_vm_group_bin_9685 (RW)
0x89: frame_vm_group_bin_2524 (RW)
0x8: frame_vm_group_bin_18295 (RW)
0x8a: frame_vm_group_bin_18601 (RW)
0x8b: frame_vm_group_bin_11537 (RW)
0x8c: frame_vm_group_bin_4355 (RW)
0x8d: frame_vm_group_bin_20451 (RW)
0x8e: frame_vm_group_bin_13254 (RW)
0x8f: frame_vm_group_bin_6082 (RW)
0x90: frame_vm_group_bin_22262 (RW)
0x91: frame_vm_group_bin_1764 (RW)
0x92: frame_vm_group_bin_7896 (RW)
0x93: frame_vm_group_bin_0732 (RW)
0x94: frame_vm_group_bin_16926 (RW)
0x95: frame_vm_group_bin_9718 (RW)
0x96: frame_vm_group_bin_2557 (RW)
0x97: frame_vm_group_bin_18634 (RW)
0x98: frame_vm_group_bin_11567 (RW)
0x99: frame_vm_group_bin_4388 (RW)
0x9: frame_vm_group_bin_11207 (RW)
0x9a: frame_vm_group_bin_20485 (RW)
0x9b: frame_vm_group_bin_13288 (RW)
0x9c: frame_vm_group_bin_6113 (RW)
0x9d: frame_vm_group_bin_22295 (RW)
0x9e: frame_vm_group_bin_15121 (RW)
0x9f: frame_vm_group_bin_7931 (RW)
0xa0: frame_vm_group_bin_0766 (RW)
0xa1: frame_vm_group_bin_16960 (RW)
0xa2: frame_vm_group_bin_9752 (RW)
0xa3: frame_vm_group_bin_2591 (RW)
0xa4: frame_vm_group_bin_18667 (RW)
0xa5: frame_vm_group_bin_19685 (RW)
0xa6: frame_vm_group_bin_4422 (RW)
0xa7: frame_vm_group_bin_20518 (RW)
0xa8: frame_vm_group_bin_13320 (RW)
0xa9: frame_vm_group_bin_6145 (RW)
0xa: frame_vm_group_bin_4022 (RW)
0xaa: frame_vm_group_bin_22328 (RW)
0xab: frame_vm_group_bin_15144 (RW)
0xac: frame_vm_group_bin_7964 (RW)
0xad: frame_vm_group_bin_0799 (RW)
0xae: frame_vm_group_bin_16993 (RW)
0xaf: frame_vm_group_bin_9785 (RW)
0xb0: frame_vm_group_bin_2624 (RW)
0xb1: frame_vm_group_bin_18700 (RW)
0xb2: frame_vm_group_bin_1051 (RW)
0xb3: frame_vm_group_bin_4455 (RW)
0xb4: frame_vm_group_bin_20551 (RW)
0xb5: frame_vm_group_bin_13353 (RW)
0xb6: frame_vm_group_bin_6178 (RW)
0xb7: frame_vm_group_bin_22360 (RW)
0xb8: frame_vm_group_bin_15176 (RW)
0xb9: frame_vm_group_bin_7995 (RW)
0xb: frame_vm_group_bin_20118 (RW)
0xba: frame_vm_group_bin_0832 (RW)
0xbb: frame_vm_group_bin_17027 (RW)
0xbc: frame_vm_group_bin_9819 (RW)
0xbd: frame_vm_group_bin_2658 (RW)
0xbe: frame_vm_group_bin_7123 (RW)
0xbf: frame_vm_group_bin_11642 (RW)
0xc0: frame_vm_group_bin_4489 (RW)
0xc1: frame_vm_group_bin_20585 (RW)
0xc2: frame_vm_group_bin_13385 (RW)
0xc3: frame_vm_group_bin_6207 (RW)
0xc4: frame_vm_group_bin_22394 (RW)
0xc5: frame_vm_group_bin_15210 (RW)
0xc6: frame_vm_group_bin_8026 (RW)
0xc7: frame_vm_group_bin_0865 (RW)
0xc8: frame_vm_group_bin_17060 (RW)
0xc9: frame_vm_group_bin_9852 (RW)
0xc: frame_vm_group_bin_12919 (RW)
0xca: frame_vm_group_bin_2691 (RW)
0xcb: frame_vm_group_bin_18764 (RW)
0xcc: frame_vm_group_bin_10422 (RW)
0xcd: frame_vm_group_bin_4522 (RW)
0xce: frame_vm_group_bin_20618 (RW)
0xcf: frame_vm_group_bin_13418 (RW)
0xd0: frame_vm_group_bin_6235 (RW)
0xd1: frame_vm_group_bin_22426 (RW)
0xd2: frame_vm_group_bin_15244 (RW)
0xd3: frame_vm_group_bin_0348 (RW)
0xd4: frame_vm_group_bin_0898 (RW)
0xd5: frame_vm_group_bin_17093 (RW)
0xd6: frame_vm_group_bin_9885 (RW)
0xd7: frame_vm_group_bin_2724 (RW)
0xd8: frame_vm_group_bin_18797 (RW)
0xd9: frame_vm_group_bin_11689 (RW)
0xd: frame_vm_group_bin_4627 (RW)
0xda: frame_vm_group_bin_4555 (RW)
0xdb: frame_vm_group_bin_12166 (RW)
0xdc: frame_vm_group_bin_13452 (RW)
0xdd: frame_vm_group_bin_6267 (RW)
0xde: frame_vm_group_bin_22460 (RW)
0xdf: frame_vm_group_bin_18823 (RW)
0xe0: frame_vm_group_bin_8087 (RW)
0xe1: frame_vm_group_bin_0932 (RW)
0xe2: frame_vm_group_bin_17127 (RW)
0xe3: frame_vm_group_bin_9918 (RW)
0xe4: frame_vm_group_bin_2758 (RW)
0xe5: frame_vm_group_bin_18832 (RW)
0xe6: frame_vm_group_bin_11718 (RW)
0xe7: frame_vm_group_bin_4583 (RW)
0xe8: frame_vm_group_bin_20684 (RW)
0xe9: frame_vm_group_bin_13485 (RW)
0xe: frame_vm_group_bin_21955 (RW)
0xea: frame_vm_group_bin_6300 (RW)
0xeb: frame_vm_group_bin_22493 (RW)
0xec: frame_vm_group_bin_15310 (RW)
0xed: frame_vm_group_bin_8119 (RW)
0xee: frame_vm_group_bin_0965 (RW)
0xef: frame_vm_group_bin_17159 (RW)
0xf0: frame_vm_group_bin_9949 (RW)
0xf1: frame_vm_group_bin_2791 (RW)
0xf2: frame_vm_group_bin_18865 (RW)
0xf3: frame_vm_group_bin_1068 (RW)
0xf4: frame_vm_group_bin_23000 (RW)
0xf5: frame_vm_group_bin_20717 (RW)
0xf6: frame_vm_group_bin_13518 (RW)
0xf7: frame_vm_group_bin_6332 (RW)
0xf8: frame_vm_group_bin_17283 (RW)
0xf9: frame_vm_group_bin_15343 (RW)
0xf: frame_vm_group_bin_14779 (RW)
0xfa: frame_vm_group_bin_8153 (RW)
0xfb: frame_vm_group_bin_0999 (RW)
0xfc: frame_vm_group_bin_11549 (RW)
0xfd: frame_vm_group_bin_9983 (RW)
0xfe: frame_vm_group_bin_2825 (RW)
0xff: frame_vm_group_bin_18899 (RW)
}
pt_vm_group_bin_0008 {
0x0: frame_vm_group_bin_22157 (RW)
0x100: frame_vm_group_bin_4888 (RW)
0x101: frame_vm_group_bin_20981 (RW)
0x102: frame_vm_group_bin_13813 (RW)
0x103: frame_vm_group_bin_6624 (RW)
0x104: frame_vm_group_bin_22820 (RW)
0x105: frame_vm_group_bin_15637 (RW)
0x106: frame_vm_group_bin_8447 (RW)
0x107: frame_vm_group_bin_1257 (RW)
0x108: frame_vm_group_bin_17459 (RW)
0x109: frame_vm_group_bin_10280 (RW)
0x10: frame_vm_group_bin_0660 (RW)
0x10a: frame_vm_group_bin_3120 (RW)
0x10b: frame_vm_group_bin_19189 (RW)
0x10c: frame_vm_group_bin_12023 (RW)
0x10d: frame_vm_group_bin_4921 (RW)
0x10e: frame_vm_group_bin_21014 (RW)
0x10f: frame_vm_group_bin_19175 (RW)
0x110: frame_vm_group_bin_6657 (RW)
0x111: frame_vm_group_bin_22853 (RW)
0x112: frame_vm_group_bin_15670 (RW)
0x113: frame_vm_group_bin_8480 (RW)
0x114: frame_vm_group_bin_1288 (RW)
0x115: frame_vm_group_bin_17478 (RW)
0x116: frame_vm_group_bin_10313 (RW)
0x117: frame_vm_group_bin_3153 (RW)
0x118: frame_vm_group_bin_19222 (RW)
0x119: frame_vm_group_bin_4907 (RW)
0x11: frame_vm_group_bin_16856 (RW)
0x11a: frame_vm_group_bin_4953 (RW)
0x11b: frame_vm_group_bin_21049 (RW)
0x11c: frame_vm_group_bin_13872 (RW)
0x11d: frame_vm_group_bin_6691 (RW)
0x11e: frame_vm_group_bin_22887 (RW)
0x11f: frame_vm_group_bin_15704 (RW)
0x120: frame_vm_group_bin_8513 (RW)
0x121: frame_vm_group_bin_1321 (RW)
0x122: frame_vm_group_bin_17501 (RW)
0x123: frame_vm_group_bin_10347 (RW)
0x124: frame_vm_group_bin_3187 (RW)
0x125: frame_vm_group_bin_19256 (RW)
0x126: frame_vm_group_bin_12083 (RW)
0x127: frame_vm_group_bin_4984 (RW)
0x128: frame_vm_group_bin_21082 (RW)
0x129: frame_vm_group_bin_13904 (RW)
0x12: frame_vm_group_bin_9647 (RW)
0x12a: frame_vm_group_bin_6723 (RW)
0x12b: frame_vm_group_bin_22920 (RW)
0x12c: frame_vm_group_bin_15737 (RW)
0x12d: frame_vm_group_bin_8546 (RW)
0x12e: frame_vm_group_bin_1354 (RW)
0x12f: frame_vm_group_bin_17529 (RW)
0x130: frame_vm_group_bin_10380 (RW)
0x131: frame_vm_group_bin_3220 (RW)
0x132: frame_vm_group_bin_19289 (RW)
0x133: frame_vm_group_bin_12115 (RW)
0x134: frame_vm_group_bin_5017 (RW)
0x135: frame_vm_group_bin_21115 (RW)
0x136: frame_vm_group_bin_13937 (RW)
0x137: frame_vm_group_bin_6756 (RW)
0x138: frame_vm_group_bin_6985 (RW)
0x139: frame_vm_group_bin_15770 (RW)
0x13: frame_vm_group_bin_2485 (RW)
0x13a: frame_vm_group_bin_8578 (RW)
0x13b: frame_vm_group_bin_1389 (RW)
0x13c: frame_vm_group_bin_17554 (RW)
0x13d: frame_vm_group_bin_10407 (RW)
0x13e: frame_vm_group_bin_3253 (RW)
0x13f: frame_vm_group_bin_19323 (RW)
0x140: frame_vm_group_bin_12149 (RW)
0x141: frame_vm_group_bin_5051 (RW)
0x142: frame_vm_group_bin_21148 (RW)
0x143: frame_vm_group_bin_13971 (RW)
0x144: frame_vm_group_bin_6789 (RW)
0x145: frame_vm_group_bin_22986 (RW)
0x146: frame_vm_group_bin_15803 (RW)
0x147: frame_vm_group_bin_8610 (RW)
0x148: frame_vm_group_bin_1422 (RW)
0x149: frame_vm_group_bin_17575 (RW)
0x14: frame_vm_group_bin_18562 (RW)
0x14a: frame_vm_group_bin_10435 (RW)
0x14b: frame_vm_group_bin_3286 (RW)
0x14c: frame_vm_group_bin_19356 (RW)
0x14d: frame_vm_group_bin_12179 (RW)
0x14e: frame_vm_group_bin_5085 (RW)
0x14f: frame_vm_group_bin_21181 (RW)
0x150: frame_vm_group_bin_14004 (RW)
0x151: frame_vm_group_bin_6820 (RW)
0x152: frame_vm_group_bin_23018 (RW)
0x153: frame_vm_group_bin_15835 (RW)
0x154: frame_vm_group_bin_8643 (RW)
0x155: frame_vm_group_bin_1455 (RW)
0x156: frame_vm_group_bin_17598 (RW)
0x157: frame_vm_group_bin_10466 (RW)
0x158: frame_vm_group_bin_3319 (RW)
0x159: frame_vm_group_bin_19389 (RW)
0x15: frame_vm_group_bin_11498 (RW)
0x15a: frame_vm_group_bin_12209 (RW)
0x15b: frame_vm_group_bin_5119 (RW)
0x15c: frame_vm_group_bin_21215 (RW)
0x15d: frame_vm_group_bin_14038 (RW)
0x15e: frame_vm_group_bin_6849 (RW)
0x15f: frame_vm_group_bin_23052 (RW)
0x160: frame_vm_group_bin_15869 (RW)
0x161: frame_vm_group_bin_8679 (RW)
0x162: frame_vm_group_bin_1489 (RW)
0x163: frame_vm_group_bin_17629 (RW)
0x164: frame_vm_group_bin_10500 (RW)
0x165: frame_vm_group_bin_3353 (RW)
0x166: frame_vm_group_bin_19422 (RW)
0x167: frame_vm_group_bin_12241 (RW)
0x168: frame_vm_group_bin_5152 (RW)
0x169: frame_vm_group_bin_21248 (RW)
0x16: frame_vm_group_bin_4314 (RW)
0x16a: frame_vm_group_bin_14071 (RW)
0x16b: frame_vm_group_bin_3845 (RW)
0x16c: frame_vm_group_bin_23085 (RW)
0x16d: frame_vm_group_bin_15902 (RW)
0x16e: frame_vm_group_bin_8711 (RW)
0x16f: frame_vm_group_bin_1522 (RW)
0x170: frame_vm_group_bin_17662 (RW)
0x171: frame_vm_group_bin_10532 (RW)
0x172: frame_vm_group_bin_3384 (RW)
0x173: frame_vm_group_bin_19453 (RW)
0x174: frame_vm_group_bin_12274 (RW)
0x175: frame_vm_group_bin_5185 (RW)
0x176: frame_vm_group_bin_21281 (RW)
0x177: frame_vm_group_bin_14104 (RW)
0x178: frame_vm_group_bin_6898 (RW)
0x179: frame_vm_group_bin_23118 (RW)
0x17: frame_vm_group_bin_20412 (RW)
0x17a: frame_vm_group_bin_15936 (RW)
0x17b: frame_vm_group_bin_8745 (RW)
0x17c: frame_vm_group_bin_1556 (RW)
0x17d: frame_vm_group_bin_17692 (RW)
0x17e: frame_vm_group_bin_10566 (RW)
0x17f: frame_vm_group_bin_3411 (RW)
0x180: frame_vm_group_bin_19486 (RW)
0x181: frame_vm_group_bin_12308 (RW)
0x182: frame_vm_group_bin_5219 (RW)
0x183: frame_vm_group_bin_21314 (RW)
0x184: frame_vm_group_bin_14138 (RW)
0x185: frame_vm_group_bin_6928 (RW)
0x186: frame_vm_group_bin_23151 (RW)
0x187: frame_vm_group_bin_15969 (RW)
0x188: frame_vm_group_bin_8778 (RW)
0x189: frame_vm_group_bin_1589 (RW)
0x18: frame_vm_group_bin_13215 (RW)
0x18a: frame_vm_group_bin_17718 (RW)
0x18b: frame_vm_group_bin_10599 (RW)
0x18c: frame_vm_group_bin_3156 (RW)
0x18d: frame_vm_group_bin_19519 (RW)
0x18e: frame_vm_group_bin_12340 (RW)
0x18f: frame_vm_group_bin_5252 (RW)
0x190: frame_vm_group_bin_21346 (RW)
0x191: frame_vm_group_bin_14171 (RW)
0x192: frame_vm_group_bin_6958 (RW)
0x193: frame_vm_group_bin_23184 (RW)
0x194: frame_vm_group_bin_16004 (RW)
0x195: frame_vm_group_bin_8811 (RW)
0x196: frame_vm_group_bin_1622 (RW)
0x197: frame_vm_group_bin_17744 (RW)
0x198: frame_vm_group_bin_10632 (RW)
0x199: frame_vm_group_bin_3458 (RW)
0x19: frame_vm_group_bin_6051 (RW)
0x19a: frame_vm_group_bin_19553 (RW)
0x19b: frame_vm_group_bin_12374 (RW)
0x19c: frame_vm_group_bin_5286 (RW)
0x19d: frame_vm_group_bin_21380 (RW)
0x19e: frame_vm_group_bin_14204 (RW)
0x19f: frame_vm_group_bin_6991 (RW)
0x1: frame_vm_group_bin_15008 (RW)
0x1a0: frame_vm_group_bin_21047 (RW)
0x1a1: frame_vm_group_bin_16038 (RW)
0x1a2: frame_vm_group_bin_8845 (RW)
0x1a3: frame_vm_group_bin_1656 (RW)
0x1a4: frame_vm_group_bin_17775 (RW)
0x1a5: frame_vm_group_bin_10664 (RW)
0x1a6: frame_vm_group_bin_12418 (RW)
0x1a7: frame_vm_group_bin_19587 (RW)
0x1a8: frame_vm_group_bin_12407 (RW)
0x1a9: frame_vm_group_bin_5318 (RW)
0x1a: frame_vm_group_bin_22224 (RW)
0x1aa: frame_vm_group_bin_21413 (RW)
0x1ab: frame_vm_group_bin_14237 (RW)
0x1ac: frame_vm_group_bin_7024 (RW)
0x1ad: frame_vm_group_bin_2421 (RW)
0x1ae: frame_vm_group_bin_16071 (RW)
0x1af: frame_vm_group_bin_8877 (RW)
0x1b0: frame_vm_group_bin_1689 (RW)
0x1b1: frame_vm_group_bin_17806 (RW)
0x1b2: frame_vm_group_bin_10697 (RW)
0x1b3: frame_vm_group_bin_3512 (RW)
0x1b4: frame_vm_group_bin_19620 (RW)
0x1b5: frame_vm_group_bin_12439 (RW)
0x1b6: frame_vm_group_bin_12765 (RW)
0x1b7: frame_vm_group_bin_21445 (RW)
0x1b8: frame_vm_group_bin_14269 (RW)
0x1b9: frame_vm_group_bin_15981 (RW)
0x1b: frame_vm_group_bin_15064 (RW)
0x1ba: frame_vm_group_bin_0004 (RW)
0x1bb: frame_vm_group_bin_16104 (RW)
0x1bc: frame_vm_group_bin_8910 (RW)
0x1bd: frame_vm_group_bin_1722 (RW)
0x1be: frame_vm_group_bin_17835 (RW)
0x1bf: frame_vm_group_bin_10730 (RW)
0x1c0: frame_vm_group_bin_3544 (RW)
0x1c1: frame_vm_group_bin_19652 (RW)
0x1c2: frame_vm_group_bin_12472 (RW)
0x1c3: frame_vm_group_bin_5382 (RW)
0x1c4: frame_vm_group_bin_21478 (RW)
0x1c5: frame_vm_group_bin_14301 (RW)
0x1c6: frame_vm_group_bin_7088 (RW)
0x1c7: frame_vm_group_bin_0021 (RW)
0x1c8: frame_vm_group_bin_16135 (RW)
0x1c9: frame_vm_group_bin_8942 (RW)
0x1c: frame_vm_group_bin_7858 (RW)
0x1ca: frame_vm_group_bin_1754 (RW)
0x1cb: frame_vm_group_bin_17862 (RW)
0x1cc: frame_vm_group_bin_10762 (RW)
0x1cd: frame_vm_group_bin_3575 (RW)
0x1ce: frame_vm_group_bin_19677 (RW)
0x1cf: frame_vm_group_bin_12504 (RW)
0x1d0: frame_vm_group_bin_5414 (RW)
0x1d1: frame_vm_group_bin_21509 (RW)
0x1d2: frame_vm_group_bin_14333 (RW)
0x1d3: frame_vm_group_bin_7119 (RW)
0x1d4: frame_vm_group_bin_0042 (RW)
0x1d5: frame_vm_group_bin_16167 (RW)
0x1d6: frame_vm_group_bin_8974 (RW)
0x1d7: frame_vm_group_bin_1786 (RW)
0x1d8: frame_vm_group_bin_17890 (RW)
0x1d9: frame_vm_group_bin_10794 (RW)
0x1d: frame_vm_group_bin_0694 (RW)
0x1da: frame_vm_group_bin_3610 (RW)
0x1db: frame_vm_group_bin_19710 (RW)
0x1dc: frame_vm_group_bin_12538 (RW)
0x1dd: frame_vm_group_bin_5448 (RW)
0x1de: frame_vm_group_bin_21543 (RW)
0x1df: frame_vm_group_bin_14367 (RW)
0x1e0: frame_vm_group_bin_7152 (RW)
0x1e1: frame_vm_group_bin_0067 (RW)
0x1e2: frame_vm_group_bin_16201 (RW)
0x1e3: frame_vm_group_bin_9008 (RW)
0x1e4: frame_vm_group_bin_1820 (RW)
0x1e5: frame_vm_group_bin_17922 (RW)
0x1e6: frame_vm_group_bin_10828 (RW)
0x1e7: frame_vm_group_bin_3643 (RW)
0x1e8: frame_vm_group_bin_19743 (RW)
0x1e9: frame_vm_group_bin_12571 (RW)
0x1e: frame_vm_group_bin_16889 (RW)
0x1ea: frame_vm_group_bin_5479 (RW)
0x1eb: frame_vm_group_bin_21576 (RW)
0x1ec: frame_vm_group_bin_14400 (RW)
0x1ed: frame_vm_group_bin_7187 (RW)
0x1ee: frame_vm_group_bin_0094 (RW)
0x1ef: frame_vm_group_bin_0997 (RW)
0x1f0: frame_vm_group_bin_9041 (RW)
0x1f1: frame_vm_group_bin_1853 (RW)
0x1f2: frame_vm_group_bin_17953 (RW)
0x1f3: frame_vm_group_bin_10861 (RW)
0x1f4: frame_vm_group_bin_3676 (RW)
0x1f5: frame_vm_group_bin_19776 (RW)
0x1f6: frame_vm_group_bin_12604 (RW)
0x1f7: frame_vm_group_bin_5512 (RW)
0x1f8: frame_vm_group_bin_21609 (RW)
0x1f9: frame_vm_group_bin_14433 (RW)
0x1f: frame_vm_group_bin_9680 (RW)
0x1fa: frame_vm_group_bin_7221 (RW)
0x1fb: frame_vm_group_bin_0120 (RW)
0x1fc: frame_vm_group_bin_16255 (RW)
0x1fd: frame_vm_group_bin_9075 (RW)
0x1fe: frame_vm_group_bin_1887 (RW)
0x1ff: frame_vm_group_bin_17985 (RW)
0x20: frame_vm_group_bin_2519 (RW)
0x21: frame_vm_group_bin_18596 (RW)
0x22: frame_vm_group_bin_11532 (RW)
0x23: frame_vm_group_bin_4350 (RW)
0x24: frame_vm_group_bin_20446 (RW)
0x25: frame_vm_group_bin_13249 (RW)
0x26: frame_vm_group_bin_6077 (RW)
0x27: frame_vm_group_bin_22257 (RW)
0x28: frame_vm_group_bin_0831 (RW)
0x29: frame_vm_group_bin_7891 (RW)
0x2: frame_vm_group_bin_7792 (RW)
0x2a: frame_vm_group_bin_0727 (RW)
0x2b: frame_vm_group_bin_16921 (RW)
0x2c: frame_vm_group_bin_9713 (RW)
0x2d: frame_vm_group_bin_2552 (RW)
0x2e: frame_vm_group_bin_18629 (RW)
0x2f: frame_vm_group_bin_11563 (RW)
0x30: frame_vm_group_bin_4383 (RW)
0x31: frame_vm_group_bin_20479 (RW)
0x32: frame_vm_group_bin_13282 (RW)
0x33: frame_vm_group_bin_6108 (RW)
0x34: frame_vm_group_bin_22289 (RW)
0x35: frame_vm_group_bin_15115 (RW)
0x36: frame_vm_group_bin_7924 (RW)
0x37: frame_vm_group_bin_0760 (RW)
0x38: frame_vm_group_bin_16954 (RW)
0x39: frame_vm_group_bin_9746 (RW)
0x3: frame_vm_group_bin_0626 (RW)
0x3a: frame_vm_group_bin_2586 (RW)
0x3b: frame_vm_group_bin_18662 (RW)
0x3c: frame_vm_group_bin_11591 (RW)
0x3d: frame_vm_group_bin_4417 (RW)
0x3e: frame_vm_group_bin_20513 (RW)
0x3f: frame_vm_group_bin_14480 (RW)
0x40: frame_vm_group_bin_6140 (RW)
0x41: frame_vm_group_bin_22323 (RW)
0x42: frame_vm_group_bin_10197 (RW)
0x43: frame_vm_group_bin_7959 (RW)
0x44: frame_vm_group_bin_0794 (RW)
0x45: frame_vm_group_bin_16988 (RW)
0x46: frame_vm_group_bin_9780 (RW)
0x47: frame_vm_group_bin_2619 (RW)
0x48: frame_vm_group_bin_18695 (RW)
0x49: frame_vm_group_bin_11616 (RW)
0x4: frame_vm_group_bin_16823 (RW)
0x4a: frame_vm_group_bin_4450 (RW)
0x4b: frame_vm_group_bin_20546 (RW)
0x4c: frame_vm_group_bin_13348 (RW)
0x4d: frame_vm_group_bin_6173 (RW)
0x4e: frame_vm_group_bin_22355 (RW)
0x4f: frame_vm_group_bin_15171 (RW)
0x50: frame_vm_group_bin_7991 (RW)
0x51: frame_vm_group_bin_0826 (RW)
0x52: frame_vm_group_bin_17021 (RW)
0x53: frame_vm_group_bin_9813 (RW)
0x54: frame_vm_group_bin_2652 (RW)
0x55: frame_vm_group_bin_18727 (RW)
0x56: frame_vm_group_bin_4834 (RW)
0x57: frame_vm_group_bin_4483 (RW)
0x58: frame_vm_group_bin_20579 (RW)
0x59: frame_vm_group_bin_13379 (RW)
0x5: frame_vm_group_bin_9614 (RW)
0x5a: frame_vm_group_bin_6205 (RW)
0x5b: frame_vm_group_bin_22389 (RW)
0x5c: frame_vm_group_bin_15205 (RW)
0x5d: frame_vm_group_bin_8022 (RW)
0x5e: frame_vm_group_bin_0860 (RW)
0x5f: frame_vm_group_bin_17055 (RW)
0x60: frame_vm_group_bin_9847 (RW)
0x61: frame_vm_group_bin_2686 (RW)
0x62: frame_vm_group_bin_18759 (RW)
0x63: frame_vm_group_bin_11661 (RW)
0x64: frame_vm_group_bin_4517 (RW)
0x65: frame_vm_group_bin_20613 (RW)
0x66: frame_vm_group_bin_13413 (RW)
0x67: frame_vm_group_bin_6231 (RW)
0x68: frame_vm_group_bin_22421 (RW)
0x69: frame_vm_group_bin_15239 (RW)
0x6: frame_vm_group_bin_2453 (RW)
0x6a: frame_vm_group_bin_8050 (RW)
0x6b: frame_vm_group_bin_0893 (RW)
0x6c: frame_vm_group_bin_17088 (RW)
0x6d: frame_vm_group_bin_9880 (RW)
0x6e: frame_vm_group_bin_2719 (RW)
0x6f: frame_vm_group_bin_18792 (RW)
0x70: frame_vm_group_bin_11685 (RW)
0x71: frame_vm_group_bin_4550 (RW)
0x72: frame_vm_group_bin_20646 (RW)
0x73: frame_vm_group_bin_13446 (RW)
0x74: frame_vm_group_bin_6262 (RW)
0x75: frame_vm_group_bin_22454 (RW)
0x76: frame_vm_group_bin_15272 (RW)
0x77: frame_vm_group_bin_8082 (RW)
0x78: frame_vm_group_bin_0926 (RW)
0x79: frame_vm_group_bin_17121 (RW)
0x7: frame_vm_group_bin_1529 (RW)
0x7a: frame_vm_group_bin_9913 (RW)
0x7b: frame_vm_group_bin_2753 (RW)
0x7c: frame_vm_group_bin_18828 (RW)
0x7d: frame_vm_group_bin_11714 (RW)
0x7e: frame_vm_group_bin_4579 (RW)
0x7f: frame_vm_group_bin_20679 (RW)
0x80: frame_vm_group_bin_13480 (RW)
0x81: frame_vm_group_bin_6295 (RW)
0x82: frame_vm_group_bin_22488 (RW)
0x83: frame_vm_group_bin_15305 (RW)
0x84: frame_vm_group_bin_8114 (RW)
0x85: frame_vm_group_bin_0960 (RW)
0x86: frame_vm_group_bin_17154 (RW)
0x87: frame_vm_group_bin_9944 (RW)
0x88: frame_vm_group_bin_2786 (RW)
0x89: frame_vm_group_bin_18860 (RW)
0x8: frame_vm_group_bin_11465 (RW)
0x8a: frame_vm_group_bin_11738 (RW)
0x8b: frame_vm_group_bin_22045 (RW)
0x8c: frame_vm_group_bin_20712 (RW)
0x8d: frame_vm_group_bin_13513 (RW)
0x8e: frame_vm_group_bin_6327 (RW)
0x8f: frame_vm_group_bin_22521 (RW)
0x90: frame_vm_group_bin_15338 (RW)
0x91: frame_vm_group_bin_8147 (RW)
0x92: frame_vm_group_bin_0993 (RW)
0x93: frame_vm_group_bin_17186 (RW)
0x94: frame_vm_group_bin_9977 (RW)
0x95: frame_vm_group_bin_2819 (RW)
0x96: frame_vm_group_bin_18893 (RW)
0x97: frame_vm_group_bin_11759 (RW)
0x98: frame_vm_group_bin_4626 (RW)
0x99: frame_vm_group_bin_20745 (RW)
0x9: frame_vm_group_bin_4281 (RW)
0x9a: frame_vm_group_bin_13547 (RW)
0x9b: frame_vm_group_bin_6361 (RW)
0x9c: frame_vm_group_bin_22554 (RW)
0x9d: frame_vm_group_bin_15372 (RW)
0x9e: frame_vm_group_bin_8181 (RW)
0x9f: frame_vm_group_bin_1024 (RW)
0xa0: frame_vm_group_bin_17218 (RW)
0xa1: frame_vm_group_bin_10011 (RW)
0xa2: frame_vm_group_bin_2853 (RW)
0xa3: frame_vm_group_bin_18927 (RW)
0xa4: frame_vm_group_bin_11785 (RW)
0xa5: frame_vm_group_bin_4658 (RW)
0xa6: frame_vm_group_bin_20779 (RW)
0xa7: frame_vm_group_bin_13580 (RW)
0xa8: frame_vm_group_bin_6391 (RW)
0xa9: frame_vm_group_bin_22587 (RW)
0xa: frame_vm_group_bin_20379 (RW)
0xaa: frame_vm_group_bin_15405 (RW)
0xab: frame_vm_group_bin_8214 (RW)
0xac: frame_vm_group_bin_1045 (RW)
0xad: frame_vm_group_bin_17250 (RW)
0xae: frame_vm_group_bin_10044 (RW)
0xaf: frame_vm_group_bin_2887 (RW)
0xb0: frame_vm_group_bin_18959 (RW)
0xb1: frame_vm_group_bin_11816 (RW)
0xb2: frame_vm_group_bin_4690 (RW)
0xb3: frame_vm_group_bin_20812 (RW)
0xb4: frame_vm_group_bin_13613 (RW)
0xb5: frame_vm_group_bin_6423 (RW)
0xb6: frame_vm_group_bin_22620 (RW)
0xb7: frame_vm_group_bin_15438 (RW)
0xb8: frame_vm_group_bin_8247 (RW)
0xb9: frame_vm_group_bin_1067 (RW)
0xb: frame_vm_group_bin_13182 (RW)
0xba: frame_vm_group_bin_17284 (RW)
0xbb: frame_vm_group_bin_10078 (RW)
0xbc: frame_vm_group_bin_2921 (RW)
0xbd: frame_vm_group_bin_18991 (RW)
0xbe: frame_vm_group_bin_11847 (RW)
0xbf: frame_vm_group_bin_4722 (RW)
0xc0: frame_vm_group_bin_20845 (RW)
0xc1: frame_vm_group_bin_13646 (RW)
0xc2: frame_vm_group_bin_6457 (RW)
0xc3: frame_vm_group_bin_22654 (RW)
0xc4: frame_vm_group_bin_15472 (RW)
0xc5: frame_vm_group_bin_8280 (RW)
0xc6: frame_vm_group_bin_1094 (RW)
0xc7: frame_vm_group_bin_17317 (RW)
0xc8: frame_vm_group_bin_10111 (RW)
0xc9: frame_vm_group_bin_2954 (RW)
0xc: frame_vm_group_bin_6025 (RW)
0xca: frame_vm_group_bin_19024 (RW)
0xcb: frame_vm_group_bin_11876 (RW)
0xcc: frame_vm_group_bin_4755 (RW)
0xcd: frame_vm_group_bin_20627 (RW)
0xce: frame_vm_group_bin_13679 (RW)
0xcf: frame_vm_group_bin_6490 (RW)
0xd0: frame_vm_group_bin_22687 (RW)
0xd1: frame_vm_group_bin_15505 (RW)
0xd2: frame_vm_group_bin_8313 (RW)
0xd3: frame_vm_group_bin_1124 (RW)
0xd4: frame_vm_group_bin_17350 (RW)
0xd5: frame_vm_group_bin_10144 (RW)
0xd6: frame_vm_group_bin_2987 (RW)
0xd7: frame_vm_group_bin_19057 (RW)
0xd8: frame_vm_group_bin_11899 (RW)
0xd9: frame_vm_group_bin_4788 (RW)
0xd: frame_vm_group_bin_22190 (RW)
0xda: frame_vm_group_bin_20897 (RW)
0xdb: frame_vm_group_bin_13712 (RW)
0xdc: frame_vm_group_bin_6524 (RW)
0xdd: frame_vm_group_bin_22721 (RW)
0xde: frame_vm_group_bin_19528 (RW)
0xdf: frame_vm_group_bin_8347 (RW)
0xe0: frame_vm_group_bin_1158 (RW)
0xe1: frame_vm_group_bin_17383 (RW)
0xe2: frame_vm_group_bin_10180 (RW)
0xe3: frame_vm_group_bin_3021 (RW)
0xe4: frame_vm_group_bin_19091 (RW)
0xe5: frame_vm_group_bin_11929 (RW)
0xe6: frame_vm_group_bin_4821 (RW)
0xe7: frame_vm_group_bin_6617 (RW)
0xe8: frame_vm_group_bin_13745 (RW)
0xe9: frame_vm_group_bin_6557 (RW)
0xe: frame_vm_group_bin_10147 (RW)
0xea: frame_vm_group_bin_22753 (RW)
0xeb: frame_vm_group_bin_15570 (RW)
0xec: frame_vm_group_bin_8380 (RW)
0xed: frame_vm_group_bin_1191 (RW)
0xee: frame_vm_group_bin_19896 (RW)
0xef: frame_vm_group_bin_10213 (RW)
0xf0: frame_vm_group_bin_3054 (RW)
0xf1: frame_vm_group_bin_19123 (RW)
0xf2: frame_vm_group_bin_11959 (RW)
0xf3: frame_vm_group_bin_4854 (RW)
0xf4: frame_vm_group_bin_11361 (RW)
0xf5: frame_vm_group_bin_13779 (RW)
0xf6: frame_vm_group_bin_6590 (RW)
0xf7: frame_vm_group_bin_22786 (RW)
0xf8: frame_vm_group_bin_15603 (RW)
0xf9: frame_vm_group_bin_8413 (RW)
0xf: frame_vm_group_bin_7825 (RW)
0xfa: frame_vm_group_bin_1225 (RW)
0xfb: frame_vm_group_bin_17436 (RW)
0xfc: frame_vm_group_bin_10247 (RW)
0xfd: frame_vm_group_bin_3088 (RW)
0xfe: frame_vm_group_bin_19156 (RW)
0xff: frame_vm_group_bin_11992 (RW)
}
pt_vm_group_bin_0010 {
0x0: frame_vm_group_bin_11626 (RW)
0x100: frame_vm_group_bin_6992 (RW)
0x101: frame_vm_group_bin_16007 (RW)
0x102: frame_vm_group_bin_16039 (RW)
0x103: frame_vm_group_bin_8846 (RW)
0x104: frame_vm_group_bin_1657 (RW)
0x105: frame_vm_group_bin_17776 (RW)
0x106: frame_vm_group_bin_10665 (RW)
0x107: frame_vm_group_bin_3486 (RW)
0x108: frame_vm_group_bin_19588 (RW)
0x109: frame_vm_group_bin_12408 (RW)
0x10: frame_vm_group_bin_2888 (RW)
0x10a: frame_vm_group_bin_5319 (RW)
0x10b: frame_vm_group_bin_21414 (RW)
0x10c: frame_vm_group_bin_14238 (RW)
0x10d: frame_vm_group_bin_7025 (RW)
0x10e: frame_vm_group_bin_23234 (RW)
0x10f: frame_vm_group_bin_16072 (RW)
0x110: frame_vm_group_bin_8878 (RW)
0x111: frame_vm_group_bin_1690 (RW)
0x112: frame_vm_group_bin_17807 (RW)
0x113: frame_vm_group_bin_10698 (RW)
0x114: frame_vm_group_bin_3513 (RW)
0x115: frame_vm_group_bin_19621 (RW)
0x116: frame_vm_group_bin_12440 (RW)
0x117: frame_vm_group_bin_5350 (RW)
0x118: frame_vm_group_bin_21446 (RW)
0x119: frame_vm_group_bin_14270 (RW)
0x11: frame_vm_group_bin_18960 (RW)
0x11a: frame_vm_group_bin_7057 (RW)
0x11b: frame_vm_group_bin_0005 (RW)
0x11c: frame_vm_group_bin_16105 (RW)
0x11d: frame_vm_group_bin_8911 (RW)
0x11e: frame_vm_group_bin_1723 (RW)
0x11f: frame_vm_group_bin_17836 (RW)
0x120: frame_vm_group_bin_10731 (RW)
0x121: frame_vm_group_bin_3545 (RW)
0x122: frame_vm_group_bin_15275 (RW)
0x123: frame_vm_group_bin_12473 (RW)
0x124: frame_vm_group_bin_5383 (RW)
0x125: frame_vm_group_bin_21479 (RW)
0x126: frame_vm_group_bin_14302 (RW)
0x127: frame_vm_group_bin_7089 (RW)
0x128: frame_vm_group_bin_0022 (RW)
0x129: frame_vm_group_bin_16136 (RW)
0x12: frame_vm_group_bin_11817 (RW)
0x12a: frame_vm_group_bin_8943 (RW)
0x12b: frame_vm_group_bin_1755 (RW)
0x12c: frame_vm_group_bin_17863 (RW)
0x12d: frame_vm_group_bin_10763 (RW)
0x12e: frame_vm_group_bin_3576 (RW)
0x12f: frame_vm_group_bin_19678 (RW)
0x130: frame_vm_group_bin_12505 (RW)
0x131: frame_vm_group_bin_5415 (RW)
0x132: frame_vm_group_bin_21510 (RW)
0x133: frame_vm_group_bin_14334 (RW)
0x134: frame_vm_group_bin_7120 (RW)
0x135: frame_vm_group_bin_0043 (RW)
0x136: frame_vm_group_bin_16168 (RW)
0x137: frame_vm_group_bin_8975 (RW)
0x138: frame_vm_group_bin_1787 (RW)
0x139: frame_vm_group_bin_17891 (RW)
0x13: frame_vm_group_bin_4691 (RW)
0x13a: frame_vm_group_bin_10796 (RW)
0x13b: frame_vm_group_bin_3611 (RW)
0x13c: frame_vm_group_bin_19711 (RW)
0x13d: frame_vm_group_bin_12539 (RW)
0x13e: frame_vm_group_bin_21753 (RW)
0x13f: frame_vm_group_bin_21544 (RW)
0x140: frame_vm_group_bin_14368 (RW)
0x141: frame_vm_group_bin_7153 (RW)
0x142: frame_vm_group_bin_0068 (RW)
0x143: frame_vm_group_bin_13000 (RW)
0x144: frame_vm_group_bin_9009 (RW)
0x145: frame_vm_group_bin_1821 (RW)
0x146: frame_vm_group_bin_17923 (RW)
0x147: frame_vm_group_bin_10829 (RW)
0x148: frame_vm_group_bin_3644 (RW)
0x149: frame_vm_group_bin_19744 (RW)
0x14: frame_vm_group_bin_20813 (RW)
0x14a: frame_vm_group_bin_12572 (RW)
0x14b: frame_vm_group_bin_5480 (RW)
0x14c: frame_vm_group_bin_21577 (RW)
0x14d: frame_vm_group_bin_14401 (RW)
0x14e: frame_vm_group_bin_7188 (RW)
0x14f: frame_vm_group_bin_0095 (RW)
0x150: frame_vm_group_bin_19200 (RW)
0x151: frame_vm_group_bin_9042 (RW)
0x152: frame_vm_group_bin_1854 (RW)
0x153: frame_vm_group_bin_17954 (RW)
0x154: frame_vm_group_bin_10862 (RW)
0x155: frame_vm_group_bin_3677 (RW)
0x156: frame_vm_group_bin_19777 (RW)
0x157: frame_vm_group_bin_12605 (RW)
0x158: frame_vm_group_bin_7736 (RW)
0x159: frame_vm_group_bin_21610 (RW)
0x15: frame_vm_group_bin_13614 (RW)
0x15a: frame_vm_group_bin_14435 (RW)
0x15b: frame_vm_group_bin_7222 (RW)
0x15c: frame_vm_group_bin_0121 (RW)
0x15d: frame_vm_group_bin_16256 (RW)
0x15e: frame_vm_group_bin_9076 (RW)
0x15f: frame_vm_group_bin_1888 (RW)
0x160: frame_vm_group_bin_17986 (RW)
0x161: frame_vm_group_bin_10896 (RW)
0x162: frame_vm_group_bin_3711 (RW)
0x163: frame_vm_group_bin_19811 (RW)
0x164: frame_vm_group_bin_12639 (RW)
0x165: frame_vm_group_bin_5546 (RW)
0x166: frame_vm_group_bin_21644 (RW)
0x167: frame_vm_group_bin_14468 (RW)
0x168: frame_vm_group_bin_7255 (RW)
0x169: frame_vm_group_bin_0142 (RW)
0x16: frame_vm_group_bin_6424 (RW)
0x16a: frame_vm_group_bin_16285 (RW)
0x16b: frame_vm_group_bin_9109 (RW)
0x16c: frame_vm_group_bin_1921 (RW)
0x16d: frame_vm_group_bin_18019 (RW)
0x16e: frame_vm_group_bin_10929 (RW)
0x16f: frame_vm_group_bin_3744 (RW)
0x170: frame_vm_group_bin_19844 (RW)
0x171: frame_vm_group_bin_18490 (RW)
0x172: frame_vm_group_bin_5579 (RW)
0x173: frame_vm_group_bin_21677 (RW)
0x174: frame_vm_group_bin_14501 (RW)
0x175: frame_vm_group_bin_7288 (RW)
0x176: frame_vm_group_bin_0164 (RW)
0x177: frame_vm_group_bin_16317 (RW)
0x178: frame_vm_group_bin_9142 (RW)
0x179: frame_vm_group_bin_1954 (RW)
0x17: frame_vm_group_bin_22621 (RW)
0x17a: frame_vm_group_bin_18053 (RW)
0x17b: frame_vm_group_bin_10963 (RW)
0x17c: frame_vm_group_bin_3778 (RW)
0x17d: frame_vm_group_bin_19878 (RW)
0x17e: frame_vm_group_bin_12692 (RW)
0x17f: frame_vm_group_bin_5612 (RW)
0x180: frame_vm_group_bin_21710 (RW)
0x181: frame_vm_group_bin_14536 (RW)
0x182: frame_vm_group_bin_7321 (RW)
0x183: frame_vm_group_bin_0195 (RW)
0x184: frame_vm_group_bin_16350 (RW)
0x185: frame_vm_group_bin_9174 (RW)
0x186: frame_vm_group_bin_1987 (RW)
0x187: frame_vm_group_bin_18084 (RW)
0x188: frame_vm_group_bin_10995 (RW)
0x189: frame_vm_group_bin_3810 (RW)
0x18: frame_vm_group_bin_15439 (RW)
0x18a: frame_vm_group_bin_19909 (RW)
0x18b: frame_vm_group_bin_12716 (RW)
0x18c: frame_vm_group_bin_5643 (RW)
0x18d: frame_vm_group_bin_21743 (RW)
0x18e: frame_vm_group_bin_14569 (RW)
0x18f: frame_vm_group_bin_7354 (RW)
0x190: frame_vm_group_bin_0226 (RW)
0x191: frame_vm_group_bin_16383 (RW)
0x192: frame_vm_group_bin_17789 (RW)
0x193: frame_vm_group_bin_2020 (RW)
0x194: frame_vm_group_bin_18116 (RW)
0x195: frame_vm_group_bin_11028 (RW)
0x196: frame_vm_group_bin_3843 (RW)
0x197: frame_vm_group_bin_19941 (RW)
0x198: frame_vm_group_bin_12741 (RW)
0x199: frame_vm_group_bin_5676 (RW)
0x19: frame_vm_group_bin_8248 (RW)
0x19a: frame_vm_group_bin_6313 (RW)
0x19b: frame_vm_group_bin_14603 (RW)
0x19c: frame_vm_group_bin_7388 (RW)
0x19d: frame_vm_group_bin_0250 (RW)
0x19e: frame_vm_group_bin_16417 (RW)
0x19f: frame_vm_group_bin_9230 (RW)
0x1: frame_vm_group_bin_17219 (RW)
0x1a0: frame_vm_group_bin_2054 (RW)
0x1a1: frame_vm_group_bin_18150 (RW)
0x1a2: frame_vm_group_bin_11062 (RW)
0x1a3: frame_vm_group_bin_3877 (RW)
0x1a4: frame_vm_group_bin_19975 (RW)
0x1a5: frame_vm_group_bin_12774 (RW)
0x1a6: frame_vm_group_bin_5710 (RW)
0x1a7: frame_vm_group_bin_21810 (RW)
0x1a8: frame_vm_group_bin_14635 (RW)
0x1a9: frame_vm_group_bin_7421 (RW)
0x1a: frame_vm_group_bin_1069 (RW)
0x1aa: frame_vm_group_bin_0273 (RW)
0x1ab: frame_vm_group_bin_16450 (RW)
0x1ac: frame_vm_group_bin_9253 (RW)
0x1ad: frame_vm_group_bin_2087 (RW)
0x1ae: frame_vm_group_bin_18183 (RW)
0x1af: frame_vm_group_bin_11095 (RW)
0x1b0: frame_vm_group_bin_3910 (RW)
0x1b1: frame_vm_group_bin_20006 (RW)
0x1b2: frame_vm_group_bin_12807 (RW)
0x1b3: frame_vm_group_bin_17167 (RW)
0x1b4: frame_vm_group_bin_21843 (RW)
0x1b5: frame_vm_group_bin_14668 (RW)
0x1b6: frame_vm_group_bin_7454 (RW)
0x1b7: frame_vm_group_bin_0302 (RW)
0x1b8: frame_vm_group_bin_16483 (RW)
0x1b9: frame_vm_group_bin_9278 (RW)
0x1b: frame_vm_group_bin_17285 (RW)
0x1ba: frame_vm_group_bin_2122 (RW)
0x1bb: frame_vm_group_bin_18216 (RW)
0x1bc: frame_vm_group_bin_11128 (RW)
0x1bd: frame_vm_group_bin_3943 (RW)
0x1be: frame_vm_group_bin_20040 (RW)
0x1bf: frame_vm_group_bin_12840 (RW)
0x1c0: frame_vm_group_bin_5766 (RW)
0x1c1: frame_vm_group_bin_21877 (RW)
0x1c2: frame_vm_group_bin_14702 (RW)
0x1c3: frame_vm_group_bin_7488 (RW)
0x1c4: frame_vm_group_bin_0334 (RW)
0x1c5: frame_vm_group_bin_16517 (RW)
0x1c6: frame_vm_group_bin_9306 (RW)
0x1c7: frame_vm_group_bin_2155 (RW)
0x1c8: frame_vm_group_bin_18249 (RW)
0x1c9: frame_vm_group_bin_11161 (RW)
0x1c: frame_vm_group_bin_10079 (RW)
0x1ca: frame_vm_group_bin_3976 (RW)
0x1cb: frame_vm_group_bin_20073 (RW)
0x1cc: frame_vm_group_bin_12873 (RW)
0x1cd: frame_vm_group_bin_5789 (RW)
0x1ce: frame_vm_group_bin_21910 (RW)
0x1cf: frame_vm_group_bin_0262 (RW)
0x1d0: frame_vm_group_bin_7520 (RW)
0x1d1: frame_vm_group_bin_0366 (RW)
0x1d2: frame_vm_group_bin_16550 (RW)
0x1d3: frame_vm_group_bin_9338 (RW)
0x1d4: frame_vm_group_bin_14503 (RW)
0x1d5: frame_vm_group_bin_18282 (RW)
0x1d6: frame_vm_group_bin_11194 (RW)
0x1d7: frame_vm_group_bin_4009 (RW)
0x1d8: frame_vm_group_bin_20106 (RW)
0x1d9: frame_vm_group_bin_12906 (RW)
0x1d: frame_vm_group_bin_2922 (RW)
0x1da: frame_vm_group_bin_5811 (RW)
0x1db: frame_vm_group_bin_21943 (RW)
0x1dc: frame_vm_group_bin_14768 (RW)
0x1dd: frame_vm_group_bin_7552 (RW)
0x1de: frame_vm_group_bin_0398 (RW)
0x1df: frame_vm_group_bin_16583 (RW)
0x1e0: frame_vm_group_bin_9372 (RW)
0x1e1: frame_vm_group_bin_2218 (RW)
0x1e2: frame_vm_group_bin_18316 (RW)
0x1e3: frame_vm_group_bin_11228 (RW)
0x1e4: frame_vm_group_bin_4043 (RW)
0x1e5: frame_vm_group_bin_20139 (RW)
0x1e6: frame_vm_group_bin_12939 (RW)
0x1e7: frame_vm_group_bin_5835 (RW)
0x1e8: frame_vm_group_bin_21976 (RW)
0x1e9: frame_vm_group_bin_14800 (RW)
0x1e: frame_vm_group_bin_18992 (RW)
0x1ea: frame_vm_group_bin_7585 (RW)
0x1eb: frame_vm_group_bin_0425 (RW)
0x1ec: frame_vm_group_bin_16615 (RW)
0x1ed: frame_vm_group_bin_9406 (RW)
0x1ee: frame_vm_group_bin_2246 (RW)
0x1ef: frame_vm_group_bin_18349 (RW)
0x1f0: frame_vm_group_bin_11261 (RW)
0x1f1: frame_vm_group_bin_4076 (RW)
0x1f2: frame_vm_group_bin_20171 (RW)
0x1f3: frame_vm_group_bin_12972 (RW)
0x1f4: frame_vm_group_bin_5859 (RW)
0x1f5: frame_vm_group_bin_22009 (RW)
0x1f6: frame_vm_group_bin_14833 (RW)
0x1f7: frame_vm_group_bin_7618 (RW)
0x1f8: frame_vm_group_bin_0458 (RW)
0x1f9: frame_vm_group_bin_16648 (RW)
0x1f: frame_vm_group_bin_11848 (RW)
0x1fa: frame_vm_group_bin_9440 (RW)
0x1fb: frame_vm_group_bin_2280 (RW)
0x1fc: frame_vm_group_bin_18383 (RW)
0x1fd: frame_vm_group_bin_11295 (RW)
0x1fe: frame_vm_group_bin_4109 (RW)
0x1ff: frame_vm_group_bin_20204 (RW)
0x20: frame_vm_group_bin_4723 (RW)
0x21: frame_vm_group_bin_10914 (RW)
0x22: frame_vm_group_bin_13647 (RW)
0x23: frame_vm_group_bin_6458 (RW)
0x24: frame_vm_group_bin_22655 (RW)
0x25: frame_vm_group_bin_15473 (RW)
0x26: frame_vm_group_bin_8281 (RW)
0x27: frame_vm_group_bin_1095 (RW)
0x28: frame_vm_group_bin_17318 (RW)
0x29: frame_vm_group_bin_10112 (RW)
0x2: frame_vm_group_bin_10012 (RW)
0x2a: frame_vm_group_bin_2955 (RW)
0x2b: frame_vm_group_bin_19025 (RW)
0x2c: frame_vm_group_bin_11877 (RW)
0x2d: frame_vm_group_bin_4756 (RW)
0x2e: frame_vm_group_bin_15556 (RW)
0x2f: frame_vm_group_bin_13680 (RW)
0x30: frame_vm_group_bin_6491 (RW)
0x31: frame_vm_group_bin_22688 (RW)
0x32: frame_vm_group_bin_15506 (RW)
0x33: frame_vm_group_bin_8314 (RW)
0x34: frame_vm_group_bin_1125 (RW)
0x35: frame_vm_group_bin_17351 (RW)
0x36: frame_vm_group_bin_10145 (RW)
0x37: frame_vm_group_bin_2988 (RW)
0x38: frame_vm_group_bin_19058 (RW)
0x39: frame_vm_group_bin_11900 (RW)
0x3: frame_vm_group_bin_2854 (RW)
0x3a: frame_vm_group_bin_4790 (RW)
0x3b: frame_vm_group_bin_20898 (RW)
0x3c: frame_vm_group_bin_13713 (RW)
0x3d: frame_vm_group_bin_6525 (RW)
0x3e: frame_vm_group_bin_22722 (RW)
0x3f: frame_vm_group_bin_15538 (RW)
0x40: frame_vm_group_bin_8348 (RW)
0x41: frame_vm_group_bin_1159 (RW)
0x42: frame_vm_group_bin_17384 (RW)
0x43: frame_vm_group_bin_10181 (RW)
0x44: frame_vm_group_bin_3022 (RW)
0x45: frame_vm_group_bin_19092 (RW)
0x46: frame_vm_group_bin_11930 (RW)
0x47: frame_vm_group_bin_4822 (RW)
0x48: frame_vm_group_bin_20923 (RW)
0x49: frame_vm_group_bin_13746 (RW)
0x4: frame_vm_group_bin_18928 (RW)
0x4a: frame_vm_group_bin_6558 (RW)
0x4b: frame_vm_group_bin_22754 (RW)
0x4c: frame_vm_group_bin_15571 (RW)
0x4d: frame_vm_group_bin_8381 (RW)
0x4e: frame_vm_group_bin_1192 (RW)
0x4f: frame_vm_group_bin_14860 (RW)
0x50: frame_vm_group_bin_10214 (RW)
0x51: frame_vm_group_bin_3055 (RW)
0x52: frame_vm_group_bin_19124 (RW)
0x53: frame_vm_group_bin_11960 (RW)
0x54: frame_vm_group_bin_4855 (RW)
0x55: frame_vm_group_bin_20950 (RW)
0x56: frame_vm_group_bin_13780 (RW)
0x57: frame_vm_group_bin_6591 (RW)
0x58: frame_vm_group_bin_22787 (RW)
0x59: frame_vm_group_bin_15604 (RW)
0x5: frame_vm_group_bin_11786 (RW)
0x5a: frame_vm_group_bin_8415 (RW)
0x5b: frame_vm_group_bin_1226 (RW)
0x5c: frame_vm_group_bin_17437 (RW)
0x5d: frame_vm_group_bin_10248 (RW)
0x5e: frame_vm_group_bin_3089 (RW)
0x5f: frame_vm_group_bin_19157 (RW)
0x60: frame_vm_group_bin_11993 (RW)
0x61: frame_vm_group_bin_4889 (RW)
0x62: frame_vm_group_bin_20982 (RW)
0x63: frame_vm_group_bin_13814 (RW)
0x64: frame_vm_group_bin_6625 (RW)
0x65: frame_vm_group_bin_22821 (RW)
0x66: frame_vm_group_bin_15638 (RW)
0x67: frame_vm_group_bin_8448 (RW)
0x68: frame_vm_group_bin_1258 (RW)
0x69: frame_vm_group_bin_0855 (RW)
0x6: frame_vm_group_bin_4659 (RW)
0x6a: frame_vm_group_bin_10281 (RW)
0x6b: frame_vm_group_bin_3121 (RW)
0x6c: frame_vm_group_bin_19190 (RW)
0x6d: frame_vm_group_bin_12024 (RW)
0x6e: frame_vm_group_bin_4922 (RW)
0x6f: frame_vm_group_bin_21015 (RW)
0x70: frame_vm_group_bin_13842 (RW)
0x71: frame_vm_group_bin_6658 (RW)
0x72: frame_vm_group_bin_22854 (RW)
0x73: frame_vm_group_bin_15671 (RW)
0x74: frame_vm_group_bin_8481 (RW)
0x75: frame_vm_group_bin_1289 (RW)
0x76: frame_vm_group_bin_17479 (RW)
0x77: frame_vm_group_bin_10314 (RW)
0x78: frame_vm_group_bin_3154 (RW)
0x79: frame_vm_group_bin_19223 (RW)
0x7: frame_vm_group_bin_20780 (RW)
0x7a: frame_vm_group_bin_12053 (RW)
0x7b: frame_vm_group_bin_4954 (RW)
0x7c: frame_vm_group_bin_21050 (RW)
0x7d: frame_vm_group_bin_13873 (RW)
0x7e: frame_vm_group_bin_6692 (RW)
0x7f: frame_vm_group_bin_22888 (RW)
0x80: frame_vm_group_bin_15705 (RW)
0x81: frame_vm_group_bin_8514 (RW)
0x82: frame_vm_group_bin_1322 (RW)
0x83: frame_vm_group_bin_17502 (RW)
0x84: frame_vm_group_bin_10348 (RW)
0x85: frame_vm_group_bin_3188 (RW)
0x86: frame_vm_group_bin_19257 (RW)
0x87: frame_vm_group_bin_12084 (RW)
0x88: frame_vm_group_bin_4985 (RW)
0x89: frame_vm_group_bin_21083 (RW)
0x8: frame_vm_group_bin_13581 (RW)
0x8a: frame_vm_group_bin_13905 (RW)
0x8b: frame_vm_group_bin_6724 (RW)
0x8c: frame_vm_group_bin_22921 (RW)
0x8d: frame_vm_group_bin_15738 (RW)
0x8e: frame_vm_group_bin_17708 (RW)
0x8f: frame_vm_group_bin_1355 (RW)
0x90: frame_vm_group_bin_17530 (RW)
0x91: frame_vm_group_bin_13403 (RW)
0x92: frame_vm_group_bin_3221 (RW)
0x93: frame_vm_group_bin_19290 (RW)
0x94: frame_vm_group_bin_12116 (RW)
0x95: frame_vm_group_bin_5018 (RW)
0x96: frame_vm_group_bin_21116 (RW)
0x97: frame_vm_group_bin_13938 (RW)
0x98: frame_vm_group_bin_11625 (RW)
0x99: frame_vm_group_bin_22953 (RW)
0x9: frame_vm_group_bin_6392 (RW)
0x9a: frame_vm_group_bin_15772 (RW)
0x9b: frame_vm_group_bin_8579 (RW)
0x9c: frame_vm_group_bin_1390 (RW)
0x9d: frame_vm_group_bin_17555 (RW)
0x9e: frame_vm_group_bin_10408 (RW)
0x9f: frame_vm_group_bin_3254 (RW)
0xa0: frame_vm_group_bin_19324 (RW)
0xa1: frame_vm_group_bin_12150 (RW)
0xa2: frame_vm_group_bin_5052 (RW)
0xa3: frame_vm_group_bin_21149 (RW)
0xa4: frame_vm_group_bin_13972 (RW)
0xa5: frame_vm_group_bin_6790 (RW)
0xa6: frame_vm_group_bin_22987 (RW)
0xa7: frame_vm_group_bin_15804 (RW)
0xa8: frame_vm_group_bin_8611 (RW)
0xa9: frame_vm_group_bin_1423 (RW)
0xa: frame_vm_group_bin_22588 (RW)
0xaa: frame_vm_group_bin_17576 (RW)
0xab: frame_vm_group_bin_10436 (RW)
0xac: frame_vm_group_bin_3287 (RW)
0xad: frame_vm_group_bin_19357 (RW)
0xae: frame_vm_group_bin_12180 (RW)
0xaf: frame_vm_group_bin_5086 (RW)
0xb0: frame_vm_group_bin_21182 (RW)
0xb1: frame_vm_group_bin_14005 (RW)
0xb2: frame_vm_group_bin_12999 (RW)
0xb3: frame_vm_group_bin_23019 (RW)
0xb4: frame_vm_group_bin_15836 (RW)
0xb5: frame_vm_group_bin_8644 (RW)
0xb6: frame_vm_group_bin_1456 (RW)
0xb7: frame_vm_group_bin_17599 (RW)
0xb8: frame_vm_group_bin_10467 (RW)
0xb9: frame_vm_group_bin_3320 (RW)
0xb: frame_vm_group_bin_15406 (RW)
0xba: frame_vm_group_bin_19391 (RW)
0xbb: frame_vm_group_bin_12210 (RW)
0xbc: frame_vm_group_bin_5120 (RW)
0xbd: frame_vm_group_bin_21216 (RW)
0xbe: frame_vm_group_bin_14039 (RW)
0xbf: frame_vm_group_bin_6850 (RW)
0xc0: frame_vm_group_bin_23053 (RW)
0xc1: frame_vm_group_bin_15870 (RW)
0xc2: frame_vm_group_bin_8680 (RW)
0xc3: frame_vm_group_bin_1490 (RW)
0xc4: frame_vm_group_bin_17630 (RW)
0xc5: frame_vm_group_bin_10501 (RW)
0xc6: frame_vm_group_bin_3354 (RW)
0xc7: frame_vm_group_bin_19423 (RW)
0xc8: frame_vm_group_bin_12242 (RW)
0xc9: frame_vm_group_bin_5153 (RW)
0xc: frame_vm_group_bin_8215 (RW)
0xca: frame_vm_group_bin_21249 (RW)
0xcb: frame_vm_group_bin_14072 (RW)
0xcc: frame_vm_group_bin_6875 (RW)
0xcd: frame_vm_group_bin_23086 (RW)
0xce: frame_vm_group_bin_15903 (RW)
0xcf: frame_vm_group_bin_8712 (RW)
0xd0: frame_vm_group_bin_1523 (RW)
0xd1: frame_vm_group_bin_17663 (RW)
0xd2: frame_vm_group_bin_10533 (RW)
0xd3: frame_vm_group_bin_3385 (RW)
0xd4: frame_vm_group_bin_19454 (RW)
0xd5: frame_vm_group_bin_12275 (RW)
0xd6: frame_vm_group_bin_5186 (RW)
0xd7: frame_vm_group_bin_21282 (RW)
0xd8: frame_vm_group_bin_14105 (RW)
0xd9: frame_vm_group_bin_6899 (RW)
0xd: frame_vm_group_bin_1046 (RW)
0xda: frame_vm_group_bin_23120 (RW)
0xdb: frame_vm_group_bin_15937 (RW)
0xdc: frame_vm_group_bin_8746 (RW)
0xdd: frame_vm_group_bin_1557 (RW)
0xde: frame_vm_group_bin_17693 (RW)
0xdf: frame_vm_group_bin_10567 (RW)
0xe0: frame_vm_group_bin_3412 (RW)
0xe1: frame_vm_group_bin_19487 (RW)
0xe2: frame_vm_group_bin_12309 (RW)
0xe3: frame_vm_group_bin_5220 (RW)
0xe4: frame_vm_group_bin_21315 (RW)
0xe5: frame_vm_group_bin_14139 (RW)
0xe6: frame_vm_group_bin_6929 (RW)
0xe7: frame_vm_group_bin_23152 (RW)
0xe8: frame_vm_group_bin_15970 (RW)
0xe9: frame_vm_group_bin_8779 (RW)
0xe: frame_vm_group_bin_17251 (RW)
0xea: frame_vm_group_bin_1590 (RW)
0xeb: frame_vm_group_bin_17719 (RW)
0xec: frame_vm_group_bin_10600 (RW)
0xed: frame_vm_group_bin_3435 (RW)
0xee: frame_vm_group_bin_19520 (RW)
0xef: frame_vm_group_bin_12341 (RW)
0xf0: frame_vm_group_bin_5253 (RW)
0xf1: frame_vm_group_bin_21347 (RW)
0xf2: frame_vm_group_bin_14172 (RW)
0xf3: frame_vm_group_bin_6959 (RW)
0xf4: frame_vm_group_bin_23185 (RW)
0xf5: frame_vm_group_bin_16005 (RW)
0xf6: frame_vm_group_bin_8812 (RW)
0xf7: frame_vm_group_bin_1623 (RW)
0xf8: frame_vm_group_bin_17745 (RW)
0xf9: frame_vm_group_bin_10633 (RW)
0xf: frame_vm_group_bin_10045 (RW)
0xfa: frame_vm_group_bin_3460 (RW)
0xfb: frame_vm_group_bin_19554 (RW)
0xfc: frame_vm_group_bin_12375 (RW)
0xfd: frame_vm_group_bin_5287 (RW)
0xfe: frame_vm_group_bin_21381 (RW)
0xff: frame_vm_group_bin_14205 (RW)
}
pt_vm_group_bin_0012 {
0x0: frame_vm_group_bin_3255 (RW)
0x100: frame_vm_group_bin_9231 (RW)
0x101: frame_vm_group_bin_2055 (RW)
0x102: frame_vm_group_bin_18151 (RW)
0x103: frame_vm_group_bin_11063 (RW)
0x104: frame_vm_group_bin_3878 (RW)
0x105: frame_vm_group_bin_19976 (RW)
0x106: frame_vm_group_bin_12775 (RW)
0x107: frame_vm_group_bin_5711 (RW)
0x108: frame_vm_group_bin_21811 (RW)
0x109: frame_vm_group_bin_14636 (RW)
0x10: frame_vm_group_bin_5087 (RW)
0x10a: frame_vm_group_bin_7422 (RW)
0x10b: frame_vm_group_bin_0274 (RW)
0x10c: frame_vm_group_bin_16451 (RW)
0x10d: frame_vm_group_bin_9254 (RW)
0x10e: frame_vm_group_bin_2088 (RW)
0x10f: frame_vm_group_bin_18184 (RW)
0x110: frame_vm_group_bin_11096 (RW)
0x111: frame_vm_group_bin_3911 (RW)
0x112: frame_vm_group_bin_20007 (RW)
0x113: frame_vm_group_bin_12808 (RW)
0x114: frame_vm_group_bin_12011 (RW)
0x115: frame_vm_group_bin_21844 (RW)
0x116: frame_vm_group_bin_14669 (RW)
0x117: frame_vm_group_bin_7455 (RW)
0x118: frame_vm_group_bin_0303 (RW)
0x119: frame_vm_group_bin_16484 (RW)
0x11: frame_vm_group_bin_21183 (RW)
0x11a: frame_vm_group_bin_9280 (RW)
0x11b: frame_vm_group_bin_2123 (RW)
0x11c: frame_vm_group_bin_18217 (RW)
0x11d: frame_vm_group_bin_11129 (RW)
0x11e: frame_vm_group_bin_3944 (RW)
0x11f: frame_vm_group_bin_20041 (RW)
0x120: frame_vm_group_bin_12841 (RW)
0x121: frame_vm_group_bin_5767 (RW)
0x122: frame_vm_group_bin_21878 (RW)
0x123: frame_vm_group_bin_14703 (RW)
0x124: frame_vm_group_bin_7489 (RW)
0x125: frame_vm_group_bin_0335 (RW)
0x126: frame_vm_group_bin_16518 (RW)
0x127: frame_vm_group_bin_9307 (RW)
0x128: frame_vm_group_bin_2156 (RW)
0x129: frame_vm_group_bin_18250 (RW)
0x12: frame_vm_group_bin_14006 (RW)
0x12a: frame_vm_group_bin_11162 (RW)
0x12b: frame_vm_group_bin_3977 (RW)
0x12c: frame_vm_group_bin_20074 (RW)
0x12d: frame_vm_group_bin_12874 (RW)
0x12e: frame_vm_group_bin_5790 (RW)
0x12f: frame_vm_group_bin_21911 (RW)
0x130: frame_vm_group_bin_14735 (RW)
0x131: frame_vm_group_bin_7521 (RW)
0x132: frame_vm_group_bin_0367 (RW)
0x133: frame_vm_group_bin_16551 (RW)
0x134: frame_vm_group_bin_9339 (RW)
0x135: frame_vm_group_bin_2188 (RW)
0x136: frame_vm_group_bin_18283 (RW)
0x137: frame_vm_group_bin_11195 (RW)
0x138: frame_vm_group_bin_4010 (RW)
0x139: frame_vm_group_bin_5653 (RW)
0x13: frame_vm_group_bin_6821 (RW)
0x13a: frame_vm_group_bin_12908 (RW)
0x13b: frame_vm_group_bin_5812 (RW)
0x13c: frame_vm_group_bin_21944 (RW)
0x13d: frame_vm_group_bin_14769 (RW)
0x13e: frame_vm_group_bin_7553 (RW)
0x13f: frame_vm_group_bin_0399 (RW)
0x140: frame_vm_group_bin_16584 (RW)
0x141: frame_vm_group_bin_9373 (RW)
0x142: frame_vm_group_bin_2219 (RW)
0x143: frame_vm_group_bin_18317 (RW)
0x144: frame_vm_group_bin_11229 (RW)
0x145: frame_vm_group_bin_4044 (RW)
0x146: frame_vm_group_bin_20140 (RW)
0x147: frame_vm_group_bin_12940 (RW)
0x148: frame_vm_group_bin_5836 (RW)
0x149: frame_vm_group_bin_21977 (RW)
0x14: frame_vm_group_bin_23020 (RW)
0x14a: frame_vm_group_bin_14801 (RW)
0x14b: frame_vm_group_bin_7586 (RW)
0x14c: frame_vm_group_bin_0426 (RW)
0x14d: frame_vm_group_bin_16616 (RW)
0x14e: frame_vm_group_bin_9407 (RW)
0x14f: frame_vm_group_bin_2247 (RW)
0x150: frame_vm_group_bin_18350 (RW)
0x151: frame_vm_group_bin_11262 (RW)
0x152: frame_vm_group_bin_4077 (RW)
0x153: frame_vm_group_bin_20172 (RW)
0x154: frame_vm_group_bin_12973 (RW)
0x155: frame_vm_group_bin_5860 (RW)
0x156: frame_vm_group_bin_10656 (RW)
0x157: frame_vm_group_bin_14834 (RW)
0x158: frame_vm_group_bin_7619 (RW)
0x159: frame_vm_group_bin_0459 (RW)
0x15: frame_vm_group_bin_15837 (RW)
0x15a: frame_vm_group_bin_16650 (RW)
0x15b: frame_vm_group_bin_9441 (RW)
0x15c: frame_vm_group_bin_2281 (RW)
0x15d: frame_vm_group_bin_18384 (RW)
0x15e: frame_vm_group_bin_11296 (RW)
0x15f: frame_vm_group_bin_4110 (RW)
0x160: frame_vm_group_bin_20205 (RW)
0x161: frame_vm_group_bin_13009 (RW)
0x162: frame_vm_group_bin_5886 (RW)
0x163: frame_vm_group_bin_22036 (RW)
0x164: frame_vm_group_bin_14868 (RW)
0x165: frame_vm_group_bin_7653 (RW)
0x166: frame_vm_group_bin_0492 (RW)
0x167: frame_vm_group_bin_16683 (RW)
0x168: frame_vm_group_bin_9474 (RW)
0x169: frame_vm_group_bin_2314 (RW)
0x16: frame_vm_group_bin_8645 (RW)
0x16a: frame_vm_group_bin_18415 (RW)
0x16b: frame_vm_group_bin_11329 (RW)
0x16c: frame_vm_group_bin_4143 (RW)
0x16d: frame_vm_group_bin_20238 (RW)
0x16e: frame_vm_group_bin_13042 (RW)
0x16f: frame_vm_group_bin_5912 (RW)
0x170: frame_vm_group_bin_22057 (RW)
0x171: frame_vm_group_bin_14901 (RW)
0x172: frame_vm_group_bin_7686 (RW)
0x173: frame_vm_group_bin_0525 (RW)
0x174: frame_vm_group_bin_16715 (RW)
0x175: frame_vm_group_bin_9507 (RW)
0x176: frame_vm_group_bin_2347 (RW)
0x177: frame_vm_group_bin_18448 (RW)
0x178: frame_vm_group_bin_11360 (RW)
0x179: frame_vm_group_bin_4175 (RW)
0x17: frame_vm_group_bin_1457 (RW)
0x17a: frame_vm_group_bin_20271 (RW)
0x17b: frame_vm_group_bin_13076 (RW)
0x17c: frame_vm_group_bin_2774 (RW)
0x17d: frame_vm_group_bin_22086 (RW)
0x17e: frame_vm_group_bin_14935 (RW)
0x17f: frame_vm_group_bin_7719 (RW)
0x180: frame_vm_group_bin_0557 (RW)
0x181: frame_vm_group_bin_16750 (RW)
0x182: frame_vm_group_bin_9541 (RW)
0x183: frame_vm_group_bin_2381 (RW)
0x184: frame_vm_group_bin_14601 (RW)
0x185: frame_vm_group_bin_11393 (RW)
0x186: frame_vm_group_bin_4208 (RW)
0x187: frame_vm_group_bin_20304 (RW)
0x188: frame_vm_group_bin_13109 (RW)
0x189: frame_vm_group_bin_5960 (RW)
0x18: frame_vm_group_bin_17600 (RW)
0x18a: frame_vm_group_bin_22117 (RW)
0x18b: frame_vm_group_bin_14968 (RW)
0x18c: frame_vm_group_bin_7752 (RW)
0x18d: frame_vm_group_bin_0588 (RW)
0x18e: frame_vm_group_bin_16783 (RW)
0x18f: frame_vm_group_bin_9574 (RW)
0x190: frame_vm_group_bin_2414 (RW)
0x191: frame_vm_group_bin_18504 (RW)
0x192: frame_vm_group_bin_11425 (RW)
0x193: frame_vm_group_bin_4241 (RW)
0x194: frame_vm_group_bin_20339 (RW)
0x195: frame_vm_group_bin_13142 (RW)
0x196: frame_vm_group_bin_5989 (RW)
0x197: frame_vm_group_bin_22150 (RW)
0x198: frame_vm_group_bin_15001 (RW)
0x199: frame_vm_group_bin_7785 (RW)
0x19: frame_vm_group_bin_10468 (RW)
0x19a: frame_vm_group_bin_0622 (RW)
0x19b: frame_vm_group_bin_16817 (RW)
0x19c: frame_vm_group_bin_9608 (RW)
0x19d: frame_vm_group_bin_2447 (RW)
0x19e: frame_vm_group_bin_18533 (RW)
0x19f: frame_vm_group_bin_11459 (RW)
0x1: frame_vm_group_bin_19325 (RW)
0x1a0: frame_vm_group_bin_4275 (RW)
0x1a1: frame_vm_group_bin_20373 (RW)
0x1a2: frame_vm_group_bin_13176 (RW)
0x1a3: frame_vm_group_bin_6020 (RW)
0x1a4: frame_vm_group_bin_22184 (RW)
0x1a5: frame_vm_group_bin_13869 (RW)
0x1a6: frame_vm_group_bin_7819 (RW)
0x1a7: frame_vm_group_bin_0654 (RW)
0x1a8: frame_vm_group_bin_16850 (RW)
0x1a9: frame_vm_group_bin_9641 (RW)
0x1a: frame_vm_group_bin_3322 (RW)
0x1aa: frame_vm_group_bin_2479 (RW)
0x1ab: frame_vm_group_bin_18558 (RW)
0x1ac: frame_vm_group_bin_11492 (RW)
0x1ad: frame_vm_group_bin_4308 (RW)
0x1ae: frame_vm_group_bin_20406 (RW)
0x1af: frame_vm_group_bin_13209 (RW)
0x1b0: frame_vm_group_bin_6048 (RW)
0x1b1: frame_vm_group_bin_22217 (RW)
0x1b2: frame_vm_group_bin_15058 (RW)
0x1b3: frame_vm_group_bin_7851 (RW)
0x1b4: frame_vm_group_bin_0687 (RW)
0x1b5: frame_vm_group_bin_16882 (RW)
0x1b6: frame_vm_group_bin_9674 (RW)
0x1b7: frame_vm_group_bin_2512 (RW)
0x1b8: frame_vm_group_bin_18589 (RW)
0x1b9: frame_vm_group_bin_11525 (RW)
0x1b: frame_vm_group_bin_19392 (RW)
0x1ba: frame_vm_group_bin_4344 (RW)
0x1bb: frame_vm_group_bin_20440 (RW)
0x1bc: frame_vm_group_bin_13243 (RW)
0x1bd: frame_vm_group_bin_6073 (RW)
0x1be: frame_vm_group_bin_22251 (RW)
0x1bf: frame_vm_group_bin_15085 (RW)
0x1c0: frame_vm_group_bin_7885 (RW)
0x1c1: frame_vm_group_bin_0721 (RW)
0x1c2: frame_vm_group_bin_16915 (RW)
0x1c3: frame_vm_group_bin_9707 (RW)
0x1c4: frame_vm_group_bin_2546 (RW)
0x1c5: frame_vm_group_bin_18623 (RW)
0x1c6: frame_vm_group_bin_13144 (RW)
0x1c7: frame_vm_group_bin_4377 (RW)
0x1c8: frame_vm_group_bin_20473 (RW)
0x1c9: frame_vm_group_bin_13276 (RW)
0x1c: frame_vm_group_bin_12211 (RW)
0x1ca: frame_vm_group_bin_6103 (RW)
0x1cb: frame_vm_group_bin_22283 (RW)
0x1cc: frame_vm_group_bin_15109 (RW)
0x1cd: frame_vm_group_bin_7918 (RW)
0x1ce: frame_vm_group_bin_0754 (RW)
0x1cf: frame_vm_group_bin_16948 (RW)
0x1d0: frame_vm_group_bin_9740 (RW)
0x1d1: frame_vm_group_bin_2579 (RW)
0x1d2: frame_vm_group_bin_18655 (RW)
0x1d3: frame_vm_group_bin_11584 (RW)
0x1d4: frame_vm_group_bin_4410 (RW)
0x1d5: frame_vm_group_bin_20506 (RW)
0x1d6: frame_vm_group_bin_13309 (RW)
0x1d7: frame_vm_group_bin_6134 (RW)
0x1d8: frame_vm_group_bin_22316 (RW)
0x1d9: frame_vm_group_bin_15135 (RW)
0x1d: frame_vm_group_bin_5121 (RW)
0x1da: frame_vm_group_bin_7953 (RW)
0x1db: frame_vm_group_bin_0788 (RW)
0x1dc: frame_vm_group_bin_16982 (RW)
0x1dd: frame_vm_group_bin_9774 (RW)
0x1de: frame_vm_group_bin_2613 (RW)
0x1df: frame_vm_group_bin_18689 (RW)
0x1e0: frame_vm_group_bin_11612 (RW)
0x1e1: frame_vm_group_bin_4444 (RW)
0x1e2: frame_vm_group_bin_20540 (RW)
0x1e3: frame_vm_group_bin_13342 (RW)
0x1e4: frame_vm_group_bin_6167 (RW)
0x1e5: frame_vm_group_bin_22349 (RW)
0x1e6: frame_vm_group_bin_15165 (RW)
0x1e7: frame_vm_group_bin_7171 (RW)
0x1e8: frame_vm_group_bin_0820 (RW)
0x1e9: frame_vm_group_bin_17015 (RW)
0x1e: frame_vm_group_bin_21217 (RW)
0x1ea: frame_vm_group_bin_9807 (RW)
0x1eb: frame_vm_group_bin_2646 (RW)
0x1ec: frame_vm_group_bin_18721 (RW)
0x1ed: frame_vm_group_bin_11634 (RW)
0x1ee: frame_vm_group_bin_4477 (RW)
0x1ef: frame_vm_group_bin_20573 (RW)
0x1f0: frame_vm_group_bin_13374 (RW)
0x1f1: frame_vm_group_bin_6198 (RW)
0x1f2: frame_vm_group_bin_22382 (RW)
0x1f3: frame_vm_group_bin_15198 (RW)
0x1f4: frame_vm_group_bin_8015 (RW)
0x1f5: frame_vm_group_bin_0853 (RW)
0x1f6: frame_vm_group_bin_17048 (RW)
0x1f7: frame_vm_group_bin_9840 (RW)
0x1f8: frame_vm_group_bin_2679 (RW)
0x1f9: frame_vm_group_bin_18752 (RW)
0x1f: frame_vm_group_bin_14040 (RW)
0x1fa: frame_vm_group_bin_11658 (RW)
0x1fb: frame_vm_group_bin_4511 (RW)
0x1fc: frame_vm_group_bin_20607 (RW)
0x1fd: frame_vm_group_bin_13407 (RW)
0x1fe: frame_vm_group_bin_6226 (RW)
0x1ff: frame_vm_group_bin_22415 (RW)
0x20: frame_vm_group_bin_6851 (RW)
0x21: frame_vm_group_bin_23054 (RW)
0x22: frame_vm_group_bin_15871 (RW)
0x23: frame_vm_group_bin_8681 (RW)
0x24: frame_vm_group_bin_1491 (RW)
0x25: frame_vm_group_bin_17631 (RW)
0x26: frame_vm_group_bin_10502 (RW)
0x27: frame_vm_group_bin_3355 (RW)
0x28: frame_vm_group_bin_19424 (RW)
0x29: frame_vm_group_bin_12243 (RW)
0x2: frame_vm_group_bin_12151 (RW)
0x2a: frame_vm_group_bin_5154 (RW)
0x2b: frame_vm_group_bin_21250 (RW)
0x2c: frame_vm_group_bin_14073 (RW)
0x2d: frame_vm_group_bin_6876 (RW)
0x2e: frame_vm_group_bin_23087 (RW)
0x2f: frame_vm_group_bin_15904 (RW)
0x30: frame_vm_group_bin_8713 (RW)
0x31: frame_vm_group_bin_1524 (RW)
0x32: frame_vm_group_bin_17664 (RW)
0x33: frame_vm_group_bin_10534 (RW)
0x34: frame_vm_group_bin_6900 (RW)
0x35: frame_vm_group_bin_5560 (RW)
0x36: frame_vm_group_bin_12276 (RW)
0x37: frame_vm_group_bin_5187 (RW)
0x38: frame_vm_group_bin_21283 (RW)
0x39: frame_vm_group_bin_14106 (RW)
0x3: frame_vm_group_bin_5053 (RW)
0x3a: frame_vm_group_bin_6901 (RW)
0x3b: frame_vm_group_bin_23121 (RW)
0x3c: frame_vm_group_bin_15938 (RW)
0x3d: frame_vm_group_bin_8747 (RW)
0x3e: frame_vm_group_bin_1558 (RW)
0x3f: frame_vm_group_bin_17694 (RW)
0x40: frame_vm_group_bin_10568 (RW)
0x41: frame_vm_group_bin_3413 (RW)
0x42: frame_vm_group_bin_19488 (RW)
0x43: frame_vm_group_bin_12310 (RW)
0x44: frame_vm_group_bin_5221 (RW)
0x45: frame_vm_group_bin_21316 (RW)
0x46: frame_vm_group_bin_14140 (RW)
0x47: frame_vm_group_bin_3037 (RW)
0x48: frame_vm_group_bin_23153 (RW)
0x49: frame_vm_group_bin_15971 (RW)
0x4: frame_vm_group_bin_21150 (RW)
0x4a: frame_vm_group_bin_8780 (RW)
0x4b: frame_vm_group_bin_1591 (RW)
0x4c: frame_vm_group_bin_17720 (RW)
0x4d: frame_vm_group_bin_10601 (RW)
0x4e: frame_vm_group_bin_16294 (RW)
0x4f: frame_vm_group_bin_19521 (RW)
0x50: frame_vm_group_bin_12342 (RW)
0x51: frame_vm_group_bin_5254 (RW)
0x52: frame_vm_group_bin_21348 (RW)
0x53: frame_vm_group_bin_14173 (RW)
0x54: frame_vm_group_bin_6960 (RW)
0x55: frame_vm_group_bin_15224 (RW)
0x56: frame_vm_group_bin_16006 (RW)
0x57: frame_vm_group_bin_8813 (RW)
0x58: frame_vm_group_bin_1624 (RW)
0x59: frame_vm_group_bin_17746 (RW)
0x5: frame_vm_group_bin_13973 (RW)
0x5a: frame_vm_group_bin_10635 (RW)
0x5b: frame_vm_group_bin_3461 (RW)
0x5c: frame_vm_group_bin_19555 (RW)
0x5d: frame_vm_group_bin_12376 (RW)
0x5e: frame_vm_group_bin_5288 (RW)
0x5f: frame_vm_group_bin_21382 (RW)
0x60: frame_vm_group_bin_14206 (RW)
0x61: frame_vm_group_bin_6993 (RW)
0x62: frame_vm_group_bin_10938 (RW)
0x63: frame_vm_group_bin_16040 (RW)
0x64: frame_vm_group_bin_8847 (RW)
0x65: frame_vm_group_bin_1658 (RW)
0x66: frame_vm_group_bin_17777 (RW)
0x67: frame_vm_group_bin_10666 (RW)
0x68: frame_vm_group_bin_3487 (RW)
0x69: frame_vm_group_bin_19589 (RW)
0x6: frame_vm_group_bin_6791 (RW)
0x6a: frame_vm_group_bin_12409 (RW)
0x6b: frame_vm_group_bin_5320 (RW)
0x6c: frame_vm_group_bin_21415 (RW)
0x6d: frame_vm_group_bin_14239 (RW)
0x6e: frame_vm_group_bin_7026 (RW)
0x6f: frame_vm_group_bin_23235 (RW)
0x70: frame_vm_group_bin_16073 (RW)
0x71: frame_vm_group_bin_8879 (RW)
0x72: frame_vm_group_bin_1691 (RW)
0x73: frame_vm_group_bin_17808 (RW)
0x74: frame_vm_group_bin_10699 (RW)
0x75: frame_vm_group_bin_3514 (RW)
0x76: frame_vm_group_bin_19622 (RW)
0x77: frame_vm_group_bin_12441 (RW)
0x78: frame_vm_group_bin_5351 (RW)
0x79: frame_vm_group_bin_21447 (RW)
0x7: frame_vm_group_bin_22988 (RW)
0x7a: frame_vm_group_bin_14272 (RW)
0x7b: frame_vm_group_bin_7058 (RW)
0x7c: frame_vm_group_bin_0006 (RW)
0x7d: frame_vm_group_bin_16106 (RW)
0x7e: frame_vm_group_bin_8912 (RW)
0x7f: frame_vm_group_bin_1724 (RW)
0x80: frame_vm_group_bin_17837 (RW)
0x81: frame_vm_group_bin_10732 (RW)
0x82: frame_vm_group_bin_3546 (RW)
0x83: frame_vm_group_bin_19653 (RW)
0x84: frame_vm_group_bin_12474 (RW)
0x85: frame_vm_group_bin_5384 (RW)
0x86: frame_vm_group_bin_21480 (RW)
0x87: frame_vm_group_bin_14303 (RW)
0x88: frame_vm_group_bin_7090 (RW)
0x89: frame_vm_group_bin_0023 (RW)
0x8: frame_vm_group_bin_15805 (RW)
0x8a: frame_vm_group_bin_16137 (RW)
0x8b: frame_vm_group_bin_8944 (RW)
0x8c: frame_vm_group_bin_1756 (RW)
0x8d: frame_vm_group_bin_17864 (RW)
0x8e: frame_vm_group_bin_10764 (RW)
0x8f: frame_vm_group_bin_3577 (RW)
0x90: frame_vm_group_bin_19679 (RW)
0x91: frame_vm_group_bin_12506 (RW)
0x92: frame_vm_group_bin_5416 (RW)
0x93: frame_vm_group_bin_21511 (RW)
0x94: frame_vm_group_bin_14335 (RW)
0x95: frame_vm_group_bin_7121 (RW)
0x96: frame_vm_group_bin_0044 (RW)
0x97: frame_vm_group_bin_16169 (RW)
0x98: frame_vm_group_bin_8976 (RW)
0x99: frame_vm_group_bin_1788 (RW)
0x9: frame_vm_group_bin_8612 (RW)
0x9a: frame_vm_group_bin_17893 (RW)
0x9b: frame_vm_group_bin_10797 (RW)
0x9c: frame_vm_group_bin_3612 (RW)
0x9d: frame_vm_group_bin_19712 (RW)
0x9e: frame_vm_group_bin_12540 (RW)
0x9f: frame_vm_group_bin_5449 (RW)
0xa0: frame_vm_group_bin_21545 (RW)
0xa1: frame_vm_group_bin_14369 (RW)
0xa2: frame_vm_group_bin_7154 (RW)
0xa3: frame_vm_group_bin_0069 (RW)
0xa4: frame_vm_group_bin_9485 (RW)
0xa5: frame_vm_group_bin_9010 (RW)
0xa6: frame_vm_group_bin_1822 (RW)
0xa7: frame_vm_group_bin_17924 (RW)
0xa8: frame_vm_group_bin_10830 (RW)
0xa9: frame_vm_group_bin_3645 (RW)
0xa: frame_vm_group_bin_1424 (RW)
0xaa: frame_vm_group_bin_19745 (RW)
0xab: frame_vm_group_bin_12573 (RW)
0xac: frame_vm_group_bin_5481 (RW)
0xad: frame_vm_group_bin_21578 (RW)
0xae: frame_vm_group_bin_14402 (RW)
0xaf: frame_vm_group_bin_7189 (RW)
0xb0: frame_vm_group_bin_0096 (RW)
0xb1: frame_vm_group_bin_16228 (RW)
0xb2: frame_vm_group_bin_9043 (RW)
0xb3: frame_vm_group_bin_1855 (RW)
0xb4: frame_vm_group_bin_17955 (RW)
0xb5: frame_vm_group_bin_10863 (RW)
0xb6: frame_vm_group_bin_3678 (RW)
0xb7: frame_vm_group_bin_19778 (RW)
0xb8: frame_vm_group_bin_12606 (RW)
0xb9: frame_vm_group_bin_5513 (RW)
0xb: frame_vm_group_bin_17577 (RW)
0xba: frame_vm_group_bin_21612 (RW)
0xbb: frame_vm_group_bin_14436 (RW)
0xbc: frame_vm_group_bin_7223 (RW)
0xbd: frame_vm_group_bin_0122 (RW)
0xbe: frame_vm_group_bin_16257 (RW)
0xbf: frame_vm_group_bin_9077 (RW)
0xc0: frame_vm_group_bin_1889 (RW)
0xc1: frame_vm_group_bin_17987 (RW)
0xc2: frame_vm_group_bin_10897 (RW)
0xc3: frame_vm_group_bin_3712 (RW)
0xc4: frame_vm_group_bin_19812 (RW)
0xc5: frame_vm_group_bin_8789 (RW)
0xc6: frame_vm_group_bin_5547 (RW)
0xc7: frame_vm_group_bin_21645 (RW)
0xc8: frame_vm_group_bin_14469 (RW)
0xc9: frame_vm_group_bin_7256 (RW)
0xc: frame_vm_group_bin_10437 (RW)
0xca: frame_vm_group_bin_0143 (RW)
0xcb: frame_vm_group_bin_16286 (RW)
0xcc: frame_vm_group_bin_9110 (RW)
0xcd: frame_vm_group_bin_1922 (RW)
0xce: frame_vm_group_bin_18020 (RW)
0xcf: frame_vm_group_bin_10930 (RW)
0xd0: frame_vm_group_bin_3745 (RW)
0xd1: frame_vm_group_bin_19845 (RW)
0xd2: frame_vm_group_bin_12667 (RW)
0xd3: frame_vm_group_bin_5580 (RW)
0xd4: frame_vm_group_bin_21678 (RW)
0xd5: frame_vm_group_bin_14502 (RW)
0xd6: frame_vm_group_bin_7289 (RW)
0xd7: frame_vm_group_bin_0165 (RW)
0xd8: frame_vm_group_bin_16318 (RW)
0xd9: frame_vm_group_bin_9143 (RW)
0xd: frame_vm_group_bin_3288 (RW)
0xda: frame_vm_group_bin_1956 (RW)
0xdb: frame_vm_group_bin_18054 (RW)
0xdc: frame_vm_group_bin_10964 (RW)
0xdd: frame_vm_group_bin_3779 (RW)
0xde: frame_vm_group_bin_19879 (RW)
0xdf: frame_vm_group_bin_12693 (RW)
0xe0: frame_vm_group_bin_16719 (RW)
0xe1: frame_vm_group_bin_21711 (RW)
0xe2: frame_vm_group_bin_14537 (RW)
0xe3: frame_vm_group_bin_7322 (RW)
0xe4: frame_vm_group_bin_0196 (RW)
0xe5: frame_vm_group_bin_16351 (RW)
0xe6: frame_vm_group_bin_9175 (RW)
0xe7: frame_vm_group_bin_1988 (RW)
0xe8: frame_vm_group_bin_18085 (RW)
0xe9: frame_vm_group_bin_10996 (RW)
0xe: frame_vm_group_bin_19358 (RW)
0xea: frame_vm_group_bin_3811 (RW)
0xeb: frame_vm_group_bin_19910 (RW)
0xec: frame_vm_group_bin_12717 (RW)
0xed: frame_vm_group_bin_5644 (RW)
0xee: frame_vm_group_bin_21744 (RW)
0xef: frame_vm_group_bin_14570 (RW)
0xf0: frame_vm_group_bin_7355 (RW)
0xf1: frame_vm_group_bin_0227 (RW)
0xf2: frame_vm_group_bin_16384 (RW)
0xf3: frame_vm_group_bin_12704 (RW)
0xf4: frame_vm_group_bin_2021 (RW)
0xf5: frame_vm_group_bin_18117 (RW)
0xf6: frame_vm_group_bin_11029 (RW)
0xf7: frame_vm_group_bin_3844 (RW)
0xf8: frame_vm_group_bin_19942 (RW)
0xf9: frame_vm_group_bin_12742 (RW)
0xf: frame_vm_group_bin_12181 (RW)
0xfa: frame_vm_group_bin_5678 (RW)
0xfb: frame_vm_group_bin_21777 (RW)
0xfc: frame_vm_group_bin_14604 (RW)
0xfd: frame_vm_group_bin_7389 (RW)
0xfe: frame_vm_group_bin_0251 (RW)
0xff: frame_vm_group_bin_16418 (RW)
}
pt_vm_group_bin_0014 {
0x0: frame_vm_group_bin_7932 (RW)
0x100: frame_vm_group_bin_13944 (RW)
0x101: frame_vm_group_bin_6762 (RW)
0x102: frame_vm_group_bin_22959 (RW)
0x103: frame_vm_group_bin_15777 (RW)
0x104: frame_vm_group_bin_8584 (RW)
0x105: frame_vm_group_bin_1395 (RW)
0x106: frame_vm_group_bin_17556 (RW)
0x107: frame_vm_group_bin_18987 (RW)
0x108: frame_vm_group_bin_3259 (RW)
0x109: frame_vm_group_bin_19329 (RW)
0x10: frame_vm_group_bin_9786 (RW)
0x10a: frame_vm_group_bin_12155 (RW)
0x10b: frame_vm_group_bin_5057 (RW)
0x10c: frame_vm_group_bin_21154 (RW)
0x10d: frame_vm_group_bin_13977 (RW)
0x10e: frame_vm_group_bin_6795 (RW)
0x10f: frame_vm_group_bin_22992 (RW)
0x110: frame_vm_group_bin_15809 (RW)
0x111: frame_vm_group_bin_8616 (RW)
0x112: frame_vm_group_bin_1428 (RW)
0x113: frame_vm_group_bin_17579 (RW)
0x114: frame_vm_group_bin_0371 (RW)
0x115: frame_vm_group_bin_3292 (RW)
0x116: frame_vm_group_bin_19362 (RW)
0x117: frame_vm_group_bin_12185 (RW)
0x118: frame_vm_group_bin_5091 (RW)
0x119: frame_vm_group_bin_21187 (RW)
0x11: frame_vm_group_bin_2625 (RW)
0x11a: frame_vm_group_bin_14011 (RW)
0x11b: frame_vm_group_bin_6826 (RW)
0x11c: frame_vm_group_bin_23025 (RW)
0x11d: frame_vm_group_bin_15842 (RW)
0x11e: frame_vm_group_bin_8650 (RW)
0x11f: frame_vm_group_bin_1462 (RW)
0x120: frame_vm_group_bin_17604 (RW)
0x121: frame_vm_group_bin_10473 (RW)
0x122: frame_vm_group_bin_3326 (RW)
0x123: frame_vm_group_bin_19396 (RW)
0x124: frame_vm_group_bin_12215 (RW)
0x125: frame_vm_group_bin_5125 (RW)
0x126: frame_vm_group_bin_21221 (RW)
0x127: frame_vm_group_bin_14044 (RW)
0x128: frame_vm_group_bin_18284 (RW)
0x129: frame_vm_group_bin_23058 (RW)
0x12: frame_vm_group_bin_18701 (RW)
0x12a: frame_vm_group_bin_15875 (RW)
0x12b: frame_vm_group_bin_8684 (RW)
0x12c: frame_vm_group_bin_1495 (RW)
0x12d: frame_vm_group_bin_17635 (RW)
0x12e: frame_vm_group_bin_10506 (RW)
0x12f: frame_vm_group_bin_3359 (RW)
0x130: frame_vm_group_bin_19428 (RW)
0x131: frame_vm_group_bin_12247 (RW)
0x132: frame_vm_group_bin_5158 (RW)
0x133: frame_vm_group_bin_21254 (RW)
0x134: frame_vm_group_bin_14077 (RW)
0x135: frame_vm_group_bin_23022 (RW)
0x136: frame_vm_group_bin_23091 (RW)
0x137: frame_vm_group_bin_15908 (RW)
0x138: frame_vm_group_bin_8717 (RW)
0x139: frame_vm_group_bin_1528 (RW)
0x13: frame_vm_group_bin_19270 (RW)
0x13a: frame_vm_group_bin_17669 (RW)
0x13b: frame_vm_group_bin_10539 (RW)
0x13c: frame_vm_group_bin_3390 (RW)
0x13d: frame_vm_group_bin_19459 (RW)
0x13e: frame_vm_group_bin_12281 (RW)
0x13f: frame_vm_group_bin_5192 (RW)
0x140: frame_vm_group_bin_21288 (RW)
0x141: frame_vm_group_bin_14111 (RW)
0x142: frame_vm_group_bin_4389 (RW)
0x143: frame_vm_group_bin_23125 (RW)
0x144: frame_vm_group_bin_15942 (RW)
0x145: frame_vm_group_bin_8751 (RW)
0x146: frame_vm_group_bin_1562 (RW)
0x147: frame_vm_group_bin_17697 (RW)
0x148: frame_vm_group_bin_10572 (RW)
0x149: frame_vm_group_bin_17601 (RW)
0x14: frame_vm_group_bin_4456 (RW)
0x14a: frame_vm_group_bin_19492 (RW)
0x14b: frame_vm_group_bin_12314 (RW)
0x14c: frame_vm_group_bin_5225 (RW)
0x14d: frame_vm_group_bin_21320 (RW)
0x14e: frame_vm_group_bin_14144 (RW)
0x14f: frame_vm_group_bin_6932 (RW)
0x150: frame_vm_group_bin_23157 (RW)
0x151: frame_vm_group_bin_15975 (RW)
0x152: frame_vm_group_bin_8784 (RW)
0x153: frame_vm_group_bin_1595 (RW)
0x154: frame_vm_group_bin_17722 (RW)
0x155: frame_vm_group_bin_10605 (RW)
0x156: frame_vm_group_bin_22292 (RW)
0x157: frame_vm_group_bin_19525 (RW)
0x158: frame_vm_group_bin_12346 (RW)
0x159: frame_vm_group_bin_5258 (RW)
0x15: frame_vm_group_bin_20552 (RW)
0x15a: frame_vm_group_bin_21353 (RW)
0x15b: frame_vm_group_bin_14178 (RW)
0x15c: frame_vm_group_bin_6965 (RW)
0x15d: frame_vm_group_bin_23190 (RW)
0x15e: frame_vm_group_bin_16011 (RW)
0x15f: frame_vm_group_bin_8818 (RW)
0x160: frame_vm_group_bin_1629 (RW)
0x161: frame_vm_group_bin_17750 (RW)
0x162: frame_vm_group_bin_10639 (RW)
0x163: frame_vm_group_bin_3655 (RW)
0x164: frame_vm_group_bin_19559 (RW)
0x165: frame_vm_group_bin_12380 (RW)
0x166: frame_vm_group_bin_5292 (RW)
0x167: frame_vm_group_bin_21386 (RW)
0x168: frame_vm_group_bin_14210 (RW)
0x169: frame_vm_group_bin_6997 (RW)
0x16: frame_vm_group_bin_13354 (RW)
0x16a: frame_vm_group_bin_23217 (RW)
0x16b: frame_vm_group_bin_16044 (RW)
0x16c: frame_vm_group_bin_8851 (RW)
0x16d: frame_vm_group_bin_1662 (RW)
0x16e: frame_vm_group_bin_17780 (RW)
0x16f: frame_vm_group_bin_10670 (RW)
0x170: frame_vm_group_bin_8294 (RW)
0x171: frame_vm_group_bin_19593 (RW)
0x172: frame_vm_group_bin_12413 (RW)
0x173: frame_vm_group_bin_5324 (RW)
0x174: frame_vm_group_bin_21419 (RW)
0x175: frame_vm_group_bin_14243 (RW)
0x176: frame_vm_group_bin_7030 (RW)
0x177: frame_vm_group_bin_21587 (RW)
0x178: frame_vm_group_bin_16077 (RW)
0x179: frame_vm_group_bin_8883 (RW)
0x17: frame_vm_group_bin_6179 (RW)
0x17a: frame_vm_group_bin_1696 (RW)
0x17b: frame_vm_group_bin_17811 (RW)
0x17c: frame_vm_group_bin_10704 (RW)
0x17d: frame_vm_group_bin_3519 (RW)
0x17e: frame_vm_group_bin_19627 (RW)
0x17f: frame_vm_group_bin_12446 (RW)
0x180: frame_vm_group_bin_5356 (RW)
0x181: frame_vm_group_bin_21452 (RW)
0x182: frame_vm_group_bin_14276 (RW)
0x183: frame_vm_group_bin_7062 (RW)
0x184: frame_vm_group_bin_0007 (RW)
0x185: frame_vm_group_bin_16110 (RW)
0x186: frame_vm_group_bin_8916 (RW)
0x187: frame_vm_group_bin_1728 (RW)
0x188: frame_vm_group_bin_17840 (RW)
0x189: frame_vm_group_bin_10736 (RW)
0x18: frame_vm_group_bin_22361 (RW)
0x18a: frame_vm_group_bin_3550 (RW)
0x18b: frame_vm_group_bin_19657 (RW)
0x18c: frame_vm_group_bin_12478 (RW)
0x18d: frame_vm_group_bin_5388 (RW)
0x18e: frame_vm_group_bin_21484 (RW)
0x18f: frame_vm_group_bin_14307 (RW)
0x190: frame_vm_group_bin_7094 (RW)
0x191: frame_vm_group_bin_0025 (RW)
0x192: frame_vm_group_bin_16141 (RW)
0x193: frame_vm_group_bin_8948 (RW)
0x194: frame_vm_group_bin_1760 (RW)
0x195: frame_vm_group_bin_17866 (RW)
0x196: frame_vm_group_bin_10769 (RW)
0x197: frame_vm_group_bin_3582 (RW)
0x198: frame_vm_group_bin_19683 (RW)
0x199: frame_vm_group_bin_12511 (RW)
0x19: frame_vm_group_bin_15177 (RW)
0x19a: frame_vm_group_bin_5422 (RW)
0x19b: frame_vm_group_bin_21517 (RW)
0x19c: frame_vm_group_bin_14341 (RW)
0x19d: frame_vm_group_bin_7127 (RW)
0x19e: frame_vm_group_bin_0048 (RW)
0x19f: frame_vm_group_bin_16175 (RW)
0x1: frame_vm_group_bin_0767 (RW)
0x1a0: frame_vm_group_bin_8982 (RW)
0x1a1: frame_vm_group_bin_1794 (RW)
0x1a2: frame_vm_group_bin_17897 (RW)
0x1a3: frame_vm_group_bin_10802 (RW)
0x1a4: frame_vm_group_bin_3617 (RW)
0x1a5: frame_vm_group_bin_19717 (RW)
0x1a6: frame_vm_group_bin_12545 (RW)
0x1a7: frame_vm_group_bin_5454 (RW)
0x1a8: frame_vm_group_bin_21550 (RW)
0x1a9: frame_vm_group_bin_14374 (RW)
0x1a: frame_vm_group_bin_7997 (RW)
0x1aa: frame_vm_group_bin_7159 (RW)
0x1ab: frame_vm_group_bin_0073 (RW)
0x1ac: frame_vm_group_bin_16206 (RW)
0x1ad: frame_vm_group_bin_9015 (RW)
0x1ae: frame_vm_group_bin_1827 (RW)
0x1af: frame_vm_group_bin_17929 (RW)
0x1b0: frame_vm_group_bin_10835 (RW)
0x1b1: frame_vm_group_bin_3650 (RW)
0x1b2: frame_vm_group_bin_19750 (RW)
0x1b3: frame_vm_group_bin_12578 (RW)
0x1b4: frame_vm_group_bin_5486 (RW)
0x1b5: frame_vm_group_bin_21583 (RW)
0x1b6: frame_vm_group_bin_14407 (RW)
0x1b7: frame_vm_group_bin_7194 (RW)
0x1b8: frame_vm_group_bin_0099 (RW)
0x1b9: frame_vm_group_bin_16233 (RW)
0x1b: frame_vm_group_bin_0833 (RW)
0x1ba: frame_vm_group_bin_9049 (RW)
0x1bb: frame_vm_group_bin_1861 (RW)
0x1bc: frame_vm_group_bin_17961 (RW)
0x1bd: frame_vm_group_bin_14434 (RW)
0x1be: frame_vm_group_bin_3684 (RW)
0x1bf: frame_vm_group_bin_19784 (RW)
0x1c0: frame_vm_group_bin_12612 (RW)
0x1c1: frame_vm_group_bin_5519 (RW)
0x1c2: frame_vm_group_bin_21617 (RW)
0x1c3: frame_vm_group_bin_14441 (RW)
0x1c4: frame_vm_group_bin_7228 (RW)
0x1c5: frame_vm_group_bin_0124 (RW)
0x1c6: frame_vm_group_bin_1506 (RW)
0x1c7: frame_vm_group_bin_9082 (RW)
0x1c8: frame_vm_group_bin_1894 (RW)
0x1c9: frame_vm_group_bin_17992 (RW)
0x1c: frame_vm_group_bin_17028 (RW)
0x1ca: frame_vm_group_bin_10902 (RW)
0x1cb: frame_vm_group_bin_3717 (RW)
0x1cc: frame_vm_group_bin_19817 (RW)
0x1cd: frame_vm_group_bin_12644 (RW)
0x1ce: frame_vm_group_bin_5552 (RW)
0x1cf: frame_vm_group_bin_21650 (RW)
0x1d0: frame_vm_group_bin_14474 (RW)
0x1d1: frame_vm_group_bin_7261 (RW)
0x1d2: frame_vm_group_bin_0145 (RW)
0x1d3: frame_vm_group_bin_16290 (RW)
0x1d4: frame_vm_group_bin_9115 (RW)
0x1d5: frame_vm_group_bin_1927 (RW)
0x1d6: frame_vm_group_bin_18025 (RW)
0x1d7: frame_vm_group_bin_10935 (RW)
0x1d8: frame_vm_group_bin_3750 (RW)
0x1d9: frame_vm_group_bin_19850 (RW)
0x1d: frame_vm_group_bin_9820 (RW)
0x1da: frame_vm_group_bin_19435 (RW)
0x1db: frame_vm_group_bin_5585 (RW)
0x1dc: frame_vm_group_bin_21683 (RW)
0x1dd: frame_vm_group_bin_14509 (RW)
0x1de: frame_vm_group_bin_7294 (RW)
0x1df: frame_vm_group_bin_0169 (RW)
0x1e0: frame_vm_group_bin_16323 (RW)
0x1e1: frame_vm_group_bin_9148 (RW)
0x1e2: frame_vm_group_bin_1960 (RW)
0x1e3: frame_vm_group_bin_18058 (RW)
0x1e4: frame_vm_group_bin_10968 (RW)
0x1e5: frame_vm_group_bin_3783 (RW)
0x1e6: frame_vm_group_bin_19883 (RW)
0x1e7: frame_vm_group_bin_0808 (RW)
0x1e8: frame_vm_group_bin_5616 (RW)
0x1e9: frame_vm_group_bin_21716 (RW)
0x1e: frame_vm_group_bin_2659 (RW)
0x1ea: frame_vm_group_bin_14542 (RW)
0x1eb: frame_vm_group_bin_7327 (RW)
0x1ec: frame_vm_group_bin_0201 (RW)
0x1ed: frame_vm_group_bin_16356 (RW)
0x1ee: frame_vm_group_bin_9180 (RW)
0x1ef: frame_vm_group_bin_1993 (RW)
0x1f0: frame_vm_group_bin_18090 (RW)
0x1f1: frame_vm_group_bin_11001 (RW)
0x1f2: frame_vm_group_bin_3816 (RW)
0x1f3: frame_vm_group_bin_19915 (RW)
0x1f4: frame_vm_group_bin_5537 (RW)
0x1f5: frame_vm_group_bin_5649 (RW)
0x1f6: frame_vm_group_bin_21749 (RW)
0x1f7: frame_vm_group_bin_14575 (RW)
0x1f8: frame_vm_group_bin_7360 (RW)
0x1f9: frame_vm_group_bin_0230 (RW)
0x1f: frame_vm_group_bin_2097 (RW)
0x1fa: frame_vm_group_bin_16390 (RW)
0x1fb: frame_vm_group_bin_9209 (RW)
0x1fc: frame_vm_group_bin_2027 (RW)
0x1fd: frame_vm_group_bin_18123 (RW)
0x1fe: frame_vm_group_bin_11035 (RW)
0x1ff: frame_vm_group_bin_3850 (RW)
0x20: frame_vm_group_bin_11643 (RW)
0x21: frame_vm_group_bin_4490 (RW)
0x22: frame_vm_group_bin_20586 (RW)
0x23: frame_vm_group_bin_13386 (RW)
0x24: frame_vm_group_bin_6208 (RW)
0x25: frame_vm_group_bin_22395 (RW)
0x26: frame_vm_group_bin_15211 (RW)
0x27: frame_vm_group_bin_13915 (RW)
0x28: frame_vm_group_bin_0866 (RW)
0x29: frame_vm_group_bin_17061 (RW)
0x2: frame_vm_group_bin_16961 (RW)
0x2a: frame_vm_group_bin_9853 (RW)
0x2b: frame_vm_group_bin_2692 (RW)
0x2c: frame_vm_group_bin_18765 (RW)
0x2d: frame_vm_group_bin_11664 (RW)
0x2e: frame_vm_group_bin_4523 (RW)
0x2f: frame_vm_group_bin_20619 (RW)
0x30: frame_vm_group_bin_13419 (RW)
0x31: frame_vm_group_bin_6236 (RW)
0x32: frame_vm_group_bin_22427 (RW)
0x33: frame_vm_group_bin_15245 (RW)
0x34: frame_vm_group_bin_8055 (RW)
0x35: frame_vm_group_bin_0899 (RW)
0x36: frame_vm_group_bin_17094 (RW)
0x37: frame_vm_group_bin_9886 (RW)
0x38: frame_vm_group_bin_2725 (RW)
0x39: frame_vm_group_bin_18798 (RW)
0x3: frame_vm_group_bin_9753 (RW)
0x3a: frame_vm_group_bin_11691 (RW)
0x3b: frame_vm_group_bin_4556 (RW)
0x3c: frame_vm_group_bin_20652 (RW)
0x3d: frame_vm_group_bin_13453 (RW)
0x3e: frame_vm_group_bin_6268 (RW)
0x3f: frame_vm_group_bin_22461 (RW)
0x40: frame_vm_group_bin_15278 (RW)
0x41: frame_vm_group_bin_8088 (RW)
0x42: frame_vm_group_bin_0933 (RW)
0x43: frame_vm_group_bin_17128 (RW)
0x44: frame_vm_group_bin_9919 (RW)
0x45: frame_vm_group_bin_2759 (RW)
0x46: frame_vm_group_bin_18833 (RW)
0x47: frame_vm_group_bin_11719 (RW)
0x48: frame_vm_group_bin_4584 (RW)
0x49: frame_vm_group_bin_20685 (RW)
0x4: frame_vm_group_bin_2592 (RW)
0x4a: frame_vm_group_bin_13486 (RW)
0x4b: frame_vm_group_bin_6301 (RW)
0x4c: frame_vm_group_bin_22494 (RW)
0x4d: frame_vm_group_bin_15311 (RW)
0x4e: frame_vm_group_bin_8120 (RW)
0x4f: frame_vm_group_bin_0966 (RW)
0x50: frame_vm_group_bin_17160 (RW)
0x51: frame_vm_group_bin_9950 (RW)
0x52: frame_vm_group_bin_2792 (RW)
0x53: frame_vm_group_bin_18866 (RW)
0x54: frame_vm_group_bin_11741 (RW)
0x55: frame_vm_group_bin_17851 (RW)
0x56: frame_vm_group_bin_20718 (RW)
0x57: frame_vm_group_bin_13519 (RW)
0x58: frame_vm_group_bin_6333 (RW)
0x59: frame_vm_group_bin_12118 (RW)
0x5: frame_vm_group_bin_18668 (RW)
0x5a: frame_vm_group_bin_15345 (RW)
0x5b: frame_vm_group_bin_8154 (RW)
0x5c: frame_vm_group_bin_1000 (RW)
0x5d: frame_vm_group_bin_6381 (RW)
0x5e: frame_vm_group_bin_9984 (RW)
0x5f: frame_vm_group_bin_2826 (RW)
0x60: frame_vm_group_bin_18900 (RW)
0x61: frame_vm_group_bin_11765 (RW)
0x62: frame_vm_group_bin_4631 (RW)
0x63: frame_vm_group_bin_20752 (RW)
0x64: frame_vm_group_bin_13553 (RW)
0x65: frame_vm_group_bin_6367 (RW)
0x66: frame_vm_group_bin_22560 (RW)
0x67: frame_vm_group_bin_15378 (RW)
0x68: frame_vm_group_bin_8187 (RW)
0x69: frame_vm_group_bin_1028 (RW)
0x6: frame_vm_group_bin_14646 (RW)
0x6a: frame_vm_group_bin_17224 (RW)
0x6b: frame_vm_group_bin_10017 (RW)
0x6c: frame_vm_group_bin_2858 (RW)
0x6d: frame_vm_group_bin_18933 (RW)
0x6e: frame_vm_group_bin_11790 (RW)
0x6f: frame_vm_group_bin_4664 (RW)
0x70: frame_vm_group_bin_20785 (RW)
0x71: frame_vm_group_bin_13586 (RW)
0x72: frame_vm_group_bin_6397 (RW)
0x73: frame_vm_group_bin_22593 (RW)
0x74: frame_vm_group_bin_15411 (RW)
0x75: frame_vm_group_bin_8220 (RW)
0x76: frame_vm_group_bin_17236 (RW)
0x77: frame_vm_group_bin_17256 (RW)
0x78: frame_vm_group_bin_10050 (RW)
0x79: frame_vm_group_bin_2893 (RW)
0x7: frame_vm_group_bin_4423 (RW)
0x7a: frame_vm_group_bin_18965 (RW)
0x7b: frame_vm_group_bin_11823 (RW)
0x7c: frame_vm_group_bin_4697 (RW)
0x7d: frame_vm_group_bin_20819 (RW)
0x7e: frame_vm_group_bin_13620 (RW)
0x7f: frame_vm_group_bin_6430 (RW)
0x80: frame_vm_group_bin_22627 (RW)
0x81: frame_vm_group_bin_15445 (RW)
0x82: frame_vm_group_bin_8254 (RW)
0x83: frame_vm_group_bin_21870 (RW)
0x84: frame_vm_group_bin_17290 (RW)
0x85: frame_vm_group_bin_10084 (RW)
0x86: frame_vm_group_bin_2927 (RW)
0x87: frame_vm_group_bin_18997 (RW)
0x88: frame_vm_group_bin_11853 (RW)
0x89: frame_vm_group_bin_4728 (RW)
0x8: frame_vm_group_bin_20519 (RW)
0x8a: frame_vm_group_bin_20849 (RW)
0x8b: frame_vm_group_bin_13652 (RW)
0x8c: frame_vm_group_bin_6463 (RW)
0x8d: frame_vm_group_bin_22660 (RW)
0x8e: frame_vm_group_bin_15478 (RW)
0x8f: frame_vm_group_bin_8286 (RW)
0x90: frame_vm_group_bin_3248 (RW)
0x91: frame_vm_group_bin_17323 (RW)
0x92: frame_vm_group_bin_10117 (RW)
0x93: frame_vm_group_bin_2960 (RW)
0x94: frame_vm_group_bin_19030 (RW)
0x95: frame_vm_group_bin_11881 (RW)
0x96: frame_vm_group_bin_4761 (RW)
0x97: frame_vm_group_bin_16508 (RW)
0x98: frame_vm_group_bin_13685 (RW)
0x99: frame_vm_group_bin_6496 (RW)
0x9: frame_vm_group_bin_13321 (RW)
0x9a: frame_vm_group_bin_22694 (RW)
0x9b: frame_vm_group_bin_10772 (RW)
0x9c: frame_vm_group_bin_8320 (RW)
0x9d: frame_vm_group_bin_1131 (RW)
0x9e: frame_vm_group_bin_17357 (RW)
0x9f: frame_vm_group_bin_10153 (RW)
0xa0: frame_vm_group_bin_2994 (RW)
0xa1: frame_vm_group_bin_19064 (RW)
0xa2: frame_vm_group_bin_11905 (RW)
0xa3: frame_vm_group_bin_4795 (RW)
0xa4: frame_vm_group_bin_21142 (RW)
0xa5: frame_vm_group_bin_13718 (RW)
0xa6: frame_vm_group_bin_6530 (RW)
0xa7: frame_vm_group_bin_22727 (RW)
0xa8: frame_vm_group_bin_15543 (RW)
0xa9: frame_vm_group_bin_8353 (RW)
0xa: frame_vm_group_bin_6146 (RW)
0xaa: frame_vm_group_bin_1164 (RW)
0xab: frame_vm_group_bin_17388 (RW)
0xac: frame_vm_group_bin_10186 (RW)
0xad: frame_vm_group_bin_3027 (RW)
0xae: frame_vm_group_bin_19097 (RW)
0xaf: frame_vm_group_bin_11935 (RW)
0xb0: frame_vm_group_bin_4827 (RW)
0xb1: frame_vm_group_bin_20928 (RW)
0xb2: frame_vm_group_bin_13751 (RW)
0xb3: frame_vm_group_bin_6563 (RW)
0xb4: frame_vm_group_bin_22759 (RW)
0xb5: frame_vm_group_bin_15576 (RW)
0xb6: frame_vm_group_bin_8386 (RW)
0xb7: frame_vm_group_bin_1197 (RW)
0xb8: frame_vm_group_bin_17414 (RW)
0xb9: frame_vm_group_bin_10219 (RW)
0xb: frame_vm_group_bin_22329 (RW)
0xba: frame_vm_group_bin_3061 (RW)
0xbb: frame_vm_group_bin_19130 (RW)
0xbc: frame_vm_group_bin_11966 (RW)
0xbd: frame_vm_group_bin_4861 (RW)
0xbe: frame_vm_group_bin_20956 (RW)
0xbf: frame_vm_group_bin_13786 (RW)
0xc0: frame_vm_group_bin_6597 (RW)
0xc1: frame_vm_group_bin_22793 (RW)
0xc2: frame_vm_group_bin_15610 (RW)
0xc3: frame_vm_group_bin_8420 (RW)
0xc4: frame_vm_group_bin_1231 (RW)
0xc5: frame_vm_group_bin_20438 (RW)
0xc6: frame_vm_group_bin_10253 (RW)
0xc7: frame_vm_group_bin_3094 (RW)
0xc8: frame_vm_group_bin_19162 (RW)
0xc9: frame_vm_group_bin_11998 (RW)
0xc: frame_vm_group_bin_6013 (RW)
0xca: frame_vm_group_bin_4894 (RW)
0xcb: frame_vm_group_bin_20987 (RW)
0xcc: frame_vm_group_bin_13818 (RW)
0xcd: frame_vm_group_bin_6630 (RW)
0xce: frame_vm_group_bin_22826 (RW)
0xcf: frame_vm_group_bin_15643 (RW)
0xd0: frame_vm_group_bin_8453 (RW)
0xd1: frame_vm_group_bin_1263 (RW)
0xd2: frame_vm_group_bin_17461 (RW)
0xd3: frame_vm_group_bin_10286 (RW)
0xd4: frame_vm_group_bin_3126 (RW)
0xd5: frame_vm_group_bin_19195 (RW)
0xd6: frame_vm_group_bin_12029 (RW)
0xd7: frame_vm_group_bin_4926 (RW)
0xd8: frame_vm_group_bin_21020 (RW)
0xd9: frame_vm_group_bin_13847 (RW)
0xd: frame_vm_group_bin_7965 (RW)
0xda: frame_vm_group_bin_6664 (RW)
0xdb: frame_vm_group_bin_22860 (RW)
0xdc: frame_vm_group_bin_15677 (RW)
0xdd: frame_vm_group_bin_8487 (RW)
0xde: frame_vm_group_bin_1295 (RW)
0xdf: frame_vm_group_bin_17482 (RW)
0xe0: frame_vm_group_bin_10320 (RW)
0xe1: frame_vm_group_bin_3160 (RW)
0xe2: frame_vm_group_bin_19229 (RW)
0xe3: frame_vm_group_bin_12057 (RW)
0xe4: frame_vm_group_bin_4958 (RW)
0xe5: frame_vm_group_bin_21055 (RW)
0xe6: frame_vm_group_bin_13877 (RW)
0xe7: frame_vm_group_bin_6697 (RW)
0xe8: frame_vm_group_bin_22893 (RW)
0xe9: frame_vm_group_bin_15710 (RW)
0xe: frame_vm_group_bin_0800 (RW)
0xea: frame_vm_group_bin_8519 (RW)
0xeb: frame_vm_group_bin_1327 (RW)
0xec: frame_vm_group_bin_17506 (RW)
0xed: frame_vm_group_bin_10353 (RW)
0xee: frame_vm_group_bin_3193 (RW)
0xef: frame_vm_group_bin_19262 (RW)
0xf0: frame_vm_group_bin_12089 (RW)
0xf1: frame_vm_group_bin_4990 (RW)
0xf2: frame_vm_group_bin_21088 (RW)
0xf3: frame_vm_group_bin_13910 (RW)
0xf4: frame_vm_group_bin_6729 (RW)
0xf5: frame_vm_group_bin_22926 (RW)
0xf6: frame_vm_group_bin_15743 (RW)
0xf7: frame_vm_group_bin_8551 (RW)
0xf8: frame_vm_group_bin_1360 (RW)
0xf9: frame_vm_group_bin_17534 (RW)
0xf: frame_vm_group_bin_16994 (RW)
0xfa: frame_vm_group_bin_10386 (RW)
0xfb: frame_vm_group_bin_3227 (RW)
0xfc: frame_vm_group_bin_19296 (RW)
0xfd: frame_vm_group_bin_12122 (RW)
0xfe: frame_vm_group_bin_5024 (RW)
0xff: frame_vm_group_bin_21122 (RW)
}
pt_vm_group_bin_0016 {
0x0: frame_vm_group_bin_10154 (RW)
0x100: frame_vm_group_bin_16176 (RW)
0x101: frame_vm_group_bin_8983 (RW)
0x102: frame_vm_group_bin_1795 (RW)
0x103: frame_vm_group_bin_17898 (RW)
0x104: frame_vm_group_bin_10803 (RW)
0x105: frame_vm_group_bin_3618 (RW)
0x106: frame_vm_group_bin_19718 (RW)
0x107: frame_vm_group_bin_12546 (RW)
0x108: frame_vm_group_bin_5455 (RW)
0x109: frame_vm_group_bin_21551 (RW)
0x10: frame_vm_group_bin_11936 (RW)
0x10a: frame_vm_group_bin_14375 (RW)
0x10b: frame_vm_group_bin_7160 (RW)
0x10c: frame_vm_group_bin_0074 (RW)
0x10d: frame_vm_group_bin_16207 (RW)
0x10e: frame_vm_group_bin_9016 (RW)
0x10f: frame_vm_group_bin_1828 (RW)
0x110: frame_vm_group_bin_17930 (RW)
0x111: frame_vm_group_bin_10836 (RW)
0x112: frame_vm_group_bin_3651 (RW)
0x113: frame_vm_group_bin_19751 (RW)
0x114: frame_vm_group_bin_12579 (RW)
0x115: frame_vm_group_bin_5487 (RW)
0x116: frame_vm_group_bin_21584 (RW)
0x117: frame_vm_group_bin_14408 (RW)
0x118: frame_vm_group_bin_7195 (RW)
0x119: frame_vm_group_bin_0100 (RW)
0x11: frame_vm_group_bin_4828 (RW)
0x11a: frame_vm_group_bin_16235 (RW)
0x11b: frame_vm_group_bin_9050 (RW)
0x11c: frame_vm_group_bin_1862 (RW)
0x11d: frame_vm_group_bin_17962 (RW)
0x11e: frame_vm_group_bin_10869 (RW)
0x11f: frame_vm_group_bin_3685 (RW)
0x120: frame_vm_group_bin_19785 (RW)
0x121: frame_vm_group_bin_12613 (RW)
0x122: frame_vm_group_bin_5520 (RW)
0x123: frame_vm_group_bin_21618 (RW)
0x124: frame_vm_group_bin_14442 (RW)
0x125: frame_vm_group_bin_7229 (RW)
0x126: frame_vm_group_bin_0125 (RW)
0x127: frame_vm_group_bin_16261 (RW)
0x128: frame_vm_group_bin_9083 (RW)
0x129: frame_vm_group_bin_1895 (RW)
0x12: frame_vm_group_bin_20929 (RW)
0x12a: frame_vm_group_bin_17993 (RW)
0x12b: frame_vm_group_bin_10903 (RW)
0x12c: frame_vm_group_bin_3718 (RW)
0x12d: frame_vm_group_bin_19818 (RW)
0x12e: frame_vm_group_bin_12645 (RW)
0x12f: frame_vm_group_bin_5553 (RW)
0x130: frame_vm_group_bin_21651 (RW)
0x131: frame_vm_group_bin_14475 (RW)
0x132: frame_vm_group_bin_7262 (RW)
0x133: frame_vm_group_bin_0146 (RW)
0x134: frame_vm_group_bin_16291 (RW)
0x135: frame_vm_group_bin_9116 (RW)
0x136: frame_vm_group_bin_1928 (RW)
0x137: frame_vm_group_bin_18026 (RW)
0x138: frame_vm_group_bin_10936 (RW)
0x139: frame_vm_group_bin_3751 (RW)
0x13: frame_vm_group_bin_13752 (RW)
0x13a: frame_vm_group_bin_19852 (RW)
0x13b: frame_vm_group_bin_12672 (RW)
0x13c: frame_vm_group_bin_5586 (RW)
0x13d: frame_vm_group_bin_21684 (RW)
0x13e: frame_vm_group_bin_14510 (RW)
0x13f: frame_vm_group_bin_7295 (RW)
0x140: frame_vm_group_bin_0170 (RW)
0x141: frame_vm_group_bin_16324 (RW)
0x142: frame_vm_group_bin_9149 (RW)
0x143: frame_vm_group_bin_1961 (RW)
0x144: frame_vm_group_bin_18059 (RW)
0x145: frame_vm_group_bin_10969 (RW)
0x146: frame_vm_group_bin_3784 (RW)
0x147: frame_vm_group_bin_19884 (RW)
0x148: frame_vm_group_bin_19010 (RW)
0x149: frame_vm_group_bin_5617 (RW)
0x14: frame_vm_group_bin_6564 (RW)
0x14a: frame_vm_group_bin_21717 (RW)
0x14b: frame_vm_group_bin_14543 (RW)
0x14c: frame_vm_group_bin_7328 (RW)
0x14d: frame_vm_group_bin_0202 (RW)
0x14e: frame_vm_group_bin_16357 (RW)
0x14f: frame_vm_group_bin_9181 (RW)
0x150: frame_vm_group_bin_1994 (RW)
0x151: frame_vm_group_bin_18091 (RW)
0x152: frame_vm_group_bin_11002 (RW)
0x153: frame_vm_group_bin_3817 (RW)
0x154: frame_vm_group_bin_19916 (RW)
0x155: frame_vm_group_bin_0393 (RW)
0x156: frame_vm_group_bin_5650 (RW)
0x157: frame_vm_group_bin_21750 (RW)
0x158: frame_vm_group_bin_14576 (RW)
0x159: frame_vm_group_bin_7361 (RW)
0x15: frame_vm_group_bin_22760 (RW)
0x15a: frame_vm_group_bin_0232 (RW)
0x15b: frame_vm_group_bin_16391 (RW)
0x15c: frame_vm_group_bin_9210 (RW)
0x15d: frame_vm_group_bin_2028 (RW)
0x15e: frame_vm_group_bin_18124 (RW)
0x15f: frame_vm_group_bin_11036 (RW)
0x160: frame_vm_group_bin_3851 (RW)
0x161: frame_vm_group_bin_19949 (RW)
0x162: frame_vm_group_bin_12748 (RW)
0x163: frame_vm_group_bin_5684 (RW)
0x164: frame_vm_group_bin_21783 (RW)
0x165: frame_vm_group_bin_14609 (RW)
0x166: frame_vm_group_bin_7395 (RW)
0x167: frame_vm_group_bin_0254 (RW)
0x168: frame_vm_group_bin_16424 (RW)
0x169: frame_vm_group_bin_18309 (RW)
0x16: frame_vm_group_bin_15577 (RW)
0x16a: frame_vm_group_bin_2061 (RW)
0x16b: frame_vm_group_bin_18157 (RW)
0x16c: frame_vm_group_bin_11069 (RW)
0x16d: frame_vm_group_bin_3884 (RW)
0x16e: frame_vm_group_bin_19982 (RW)
0x16f: frame_vm_group_bin_12781 (RW)
0x170: frame_vm_group_bin_5717 (RW)
0x171: frame_vm_group_bin_21817 (RW)
0x172: frame_vm_group_bin_14642 (RW)
0x173: frame_vm_group_bin_7428 (RW)
0x174: frame_vm_group_bin_0278 (RW)
0x175: frame_vm_group_bin_16457 (RW)
0x176: frame_vm_group_bin_23046 (RW)
0x177: frame_vm_group_bin_2094 (RW)
0x178: frame_vm_group_bin_18190 (RW)
0x179: frame_vm_group_bin_11102 (RW)
0x17: frame_vm_group_bin_8387 (RW)
0x17a: frame_vm_group_bin_3918 (RW)
0x17b: frame_vm_group_bin_20014 (RW)
0x17c: frame_vm_group_bin_12815 (RW)
0x17d: frame_vm_group_bin_12929 (RW)
0x17e: frame_vm_group_bin_21851 (RW)
0x17f: frame_vm_group_bin_14676 (RW)
0x180: frame_vm_group_bin_7462 (RW)
0x181: frame_vm_group_bin_0309 (RW)
0x182: frame_vm_group_bin_16491 (RW)
0x183: frame_vm_group_bin_4413 (RW)
0x184: frame_vm_group_bin_2129 (RW)
0x185: frame_vm_group_bin_18223 (RW)
0x186: frame_vm_group_bin_11135 (RW)
0x187: frame_vm_group_bin_3950 (RW)
0x188: frame_vm_group_bin_20047 (RW)
0x189: frame_vm_group_bin_12847 (RW)
0x18: frame_vm_group_bin_1198 (RW)
0x18a: frame_vm_group_bin_17622 (RW)
0x18b: frame_vm_group_bin_21884 (RW)
0x18c: frame_vm_group_bin_14709 (RW)
0x18d: frame_vm_group_bin_7495 (RW)
0x18e: frame_vm_group_bin_0341 (RW)
0x18f: frame_vm_group_bin_16524 (RW)
0x190: frame_vm_group_bin_9312 (RW)
0x191: frame_vm_group_bin_2162 (RW)
0x192: frame_vm_group_bin_18256 (RW)
0x193: frame_vm_group_bin_11168 (RW)
0x194: frame_vm_group_bin_3983 (RW)
0x195: frame_vm_group_bin_20080 (RW)
0x196: frame_vm_group_bin_12880 (RW)
0x197: frame_vm_group_bin_22317 (RW)
0x198: frame_vm_group_bin_20875 (RW)
0x199: frame_vm_group_bin_14741 (RW)
0x19: frame_vm_group_bin_17415 (RW)
0x19a: frame_vm_group_bin_7528 (RW)
0x19b: frame_vm_group_bin_0373 (RW)
0x19c: frame_vm_group_bin_16557 (RW)
0x19d: frame_vm_group_bin_9346 (RW)
0x19e: frame_vm_group_bin_2195 (RW)
0x19f: frame_vm_group_bin_18290 (RW)
0x1: frame_vm_group_bin_2995 (RW)
0x1a0: frame_vm_group_bin_11202 (RW)
0x1a1: frame_vm_group_bin_4017 (RW)
0x1a2: frame_vm_group_bin_20113 (RW)
0x1a3: frame_vm_group_bin_12914 (RW)
0x1a4: frame_vm_group_bin_5815 (RW)
0x1a5: frame_vm_group_bin_21950 (RW)
0x1a6: frame_vm_group_bin_14775 (RW)
0x1a7: frame_vm_group_bin_7559 (RW)
0x1a8: frame_vm_group_bin_0403 (RW)
0x1a9: frame_vm_group_bin_16590 (RW)
0x1a: frame_vm_group_bin_10221 (RW)
0x1aa: frame_vm_group_bin_9379 (RW)
0x1ab: frame_vm_group_bin_2224 (RW)
0x1ac: frame_vm_group_bin_18323 (RW)
0x1ad: frame_vm_group_bin_11235 (RW)
0x1ae: frame_vm_group_bin_4050 (RW)
0x1af: frame_vm_group_bin_20146 (RW)
0x1b0: frame_vm_group_bin_12946 (RW)
0x1b1: frame_vm_group_bin_5840 (RW)
0x1b2: frame_vm_group_bin_21983 (RW)
0x1b3: frame_vm_group_bin_14807 (RW)
0x1b4: frame_vm_group_bin_7592 (RW)
0x1b5: frame_vm_group_bin_0432 (RW)
0x1b6: frame_vm_group_bin_16622 (RW)
0x1b7: frame_vm_group_bin_9413 (RW)
0x1b8: frame_vm_group_bin_2253 (RW)
0x1b9: frame_vm_group_bin_18356 (RW)
0x1b: frame_vm_group_bin_3062 (RW)
0x1ba: frame_vm_group_bin_11269 (RW)
0x1bb: frame_vm_group_bin_4084 (RW)
0x1bc: frame_vm_group_bin_20179 (RW)
0x1bd: frame_vm_group_bin_12980 (RW)
0x1be: frame_vm_group_bin_5864 (RW)
0x1bf: frame_vm_group_bin_22016 (RW)
0x1c0: frame_vm_group_bin_14841 (RW)
0x1c1: frame_vm_group_bin_7626 (RW)
0x1c2: frame_vm_group_bin_0466 (RW)
0x1c3: frame_vm_group_bin_16656 (RW)
0x1c4: frame_vm_group_bin_9447 (RW)
0x1c5: frame_vm_group_bin_2287 (RW)
0x1c6: frame_vm_group_bin_18390 (RW)
0x1c7: frame_vm_group_bin_11302 (RW)
0x1c8: frame_vm_group_bin_4116 (RW)
0x1c9: frame_vm_group_bin_20211 (RW)
0x1c: frame_vm_group_bin_6359 (RW)
0x1ca: frame_vm_group_bin_13015 (RW)
0x1cb: frame_vm_group_bin_5890 (RW)
0x1cc: frame_vm_group_bin_16252 (RW)
0x1cd: frame_vm_group_bin_14874 (RW)
0x1ce: frame_vm_group_bin_7659 (RW)
0x1cf: frame_vm_group_bin_0498 (RW)
0x1d0: frame_vm_group_bin_16689 (RW)
0x1d1: frame_vm_group_bin_9480 (RW)
0x1d2: frame_vm_group_bin_2320 (RW)
0x1d3: frame_vm_group_bin_18421 (RW)
0x1d4: frame_vm_group_bin_11335 (RW)
0x1d5: frame_vm_group_bin_4149 (RW)
0x1d6: frame_vm_group_bin_20244 (RW)
0x1d7: frame_vm_group_bin_13048 (RW)
0x1d8: frame_vm_group_bin_5916 (RW)
0x1d9: frame_vm_group_bin_22062 (RW)
0x1d: frame_vm_group_bin_11967 (RW)
0x1da: frame_vm_group_bin_14908 (RW)
0x1db: frame_vm_group_bin_7693 (RW)
0x1dc: frame_vm_group_bin_0531 (RW)
0x1dd: frame_vm_group_bin_16723 (RW)
0x1de: frame_vm_group_bin_9514 (RW)
0x1df: frame_vm_group_bin_2354 (RW)
0x1e0: frame_vm_group_bin_18455 (RW)
0x1e1: frame_vm_group_bin_11367 (RW)
0x1e2: frame_vm_group_bin_4182 (RW)
0x1e3: frame_vm_group_bin_20277 (RW)
0x1e4: frame_vm_group_bin_13082 (RW)
0x1e5: frame_vm_group_bin_5940 (RW)
0x1e6: frame_vm_group_bin_22091 (RW)
0x1e7: frame_vm_group_bin_14941 (RW)
0x1e8: frame_vm_group_bin_7725 (RW)
0x1e9: frame_vm_group_bin_0562 (RW)
0x1e: frame_vm_group_bin_4862 (RW)
0x1ea: frame_vm_group_bin_16756 (RW)
0x1eb: frame_vm_group_bin_9547 (RW)
0x1ec: frame_vm_group_bin_2387 (RW)
0x1ed: frame_vm_group_bin_15533 (RW)
0x1ee: frame_vm_group_bin_11399 (RW)
0x1ef: frame_vm_group_bin_4214 (RW)
0x1f0: frame_vm_group_bin_20310 (RW)
0x1f1: frame_vm_group_bin_13115 (RW)
0x1f2: frame_vm_group_bin_5965 (RW)
0x1f3: frame_vm_group_bin_22123 (RW)
0x1f4: frame_vm_group_bin_14974 (RW)
0x1f5: frame_vm_group_bin_7758 (RW)
0x1f6: frame_vm_group_bin_0594 (RW)
0x1f7: frame_vm_group_bin_16789 (RW)
0x1f8: frame_vm_group_bin_9580 (RW)
0x1f9: frame_vm_group_bin_2420 (RW)
0x1f: frame_vm_group_bin_20957 (RW)
0x1fa: frame_vm_group_bin_18511 (RW)
0x1fb: frame_vm_group_bin_11432 (RW)
0x1fc: frame_vm_group_bin_4248 (RW)
0x1fd: frame_vm_group_bin_20346 (RW)
0x1fe: frame_vm_group_bin_13149 (RW)
0x1ff: frame_vm_group_bin_5994 (RW)
0x20: frame_vm_group_bin_13787 (RW)
0x21: frame_vm_group_bin_6598 (RW)
0x22: frame_vm_group_bin_22794 (RW)
0x23: frame_vm_group_bin_15611 (RW)
0x24: frame_vm_group_bin_8421 (RW)
0x25: frame_vm_group_bin_1232 (RW)
0x26: frame_vm_group_bin_15368 (RW)
0x27: frame_vm_group_bin_10254 (RW)
0x28: frame_vm_group_bin_3095 (RW)
0x29: frame_vm_group_bin_19163 (RW)
0x2: frame_vm_group_bin_19065 (RW)
0x2a: frame_vm_group_bin_11999 (RW)
0x2b: frame_vm_group_bin_4895 (RW)
0x2c: frame_vm_group_bin_20988 (RW)
0x2d: frame_vm_group_bin_13819 (RW)
0x2e: frame_vm_group_bin_6631 (RW)
0x2f: frame_vm_group_bin_22827 (RW)
0x30: frame_vm_group_bin_15644 (RW)
0x31: frame_vm_group_bin_8454 (RW)
0x32: frame_vm_group_bin_1264 (RW)
0x33: frame_vm_group_bin_17462 (RW)
0x34: frame_vm_group_bin_10287 (RW)
0x35: frame_vm_group_bin_3127 (RW)
0x36: frame_vm_group_bin_19196 (RW)
0x37: frame_vm_group_bin_14292 (RW)
0x38: frame_vm_group_bin_4927 (RW)
0x39: frame_vm_group_bin_21021 (RW)
0x3: frame_vm_group_bin_11906 (RW)
0x3a: frame_vm_group_bin_13849 (RW)
0x3b: frame_vm_group_bin_6665 (RW)
0x3c: frame_vm_group_bin_22861 (RW)
0x3d: frame_vm_group_bin_15678 (RW)
0x3e: frame_vm_group_bin_8488 (RW)
0x3f: frame_vm_group_bin_1296 (RW)
0x40: frame_vm_group_bin_17483 (RW)
0x41: frame_vm_group_bin_10321 (RW)
0x42: frame_vm_group_bin_3161 (RW)
0x43: frame_vm_group_bin_19230 (RW)
0x44: frame_vm_group_bin_12058 (RW)
0x45: frame_vm_group_bin_4959 (RW)
0x46: frame_vm_group_bin_21056 (RW)
0x47: frame_vm_group_bin_13878 (RW)
0x48: frame_vm_group_bin_6698 (RW)
0x49: frame_vm_group_bin_22894 (RW)
0x4: frame_vm_group_bin_4796 (RW)
0x4a: frame_vm_group_bin_15711 (RW)
0x4b: frame_vm_group_bin_8520 (RW)
0x4c: frame_vm_group_bin_1328 (RW)
0x4d: frame_vm_group_bin_17507 (RW)
0x4e: frame_vm_group_bin_10354 (RW)
0x4f: frame_vm_group_bin_3194 (RW)
0x50: frame_vm_group_bin_19263 (RW)
0x51: frame_vm_group_bin_12090 (RW)
0x52: frame_vm_group_bin_4991 (RW)
0x53: frame_vm_group_bin_21089 (RW)
0x54: frame_vm_group_bin_13911 (RW)
0x55: frame_vm_group_bin_6730 (RW)
0x56: frame_vm_group_bin_22927 (RW)
0x57: frame_vm_group_bin_15744 (RW)
0x58: frame_vm_group_bin_8552 (RW)
0x59: frame_vm_group_bin_1363 (RW)
0x5: frame_vm_group_bin_16102 (RW)
0x5a: frame_vm_group_bin_17536 (RW)
0x5b: frame_vm_group_bin_10387 (RW)
0x5c: frame_vm_group_bin_3228 (RW)
0x5d: frame_vm_group_bin_19297 (RW)
0x5e: frame_vm_group_bin_12123 (RW)
0x5f: frame_vm_group_bin_5025 (RW)
0x60: frame_vm_group_bin_21123 (RW)
0x61: frame_vm_group_bin_13945 (RW)
0x62: frame_vm_group_bin_6763 (RW)
0x63: frame_vm_group_bin_22960 (RW)
0x64: frame_vm_group_bin_15778 (RW)
0x65: frame_vm_group_bin_8585 (RW)
0x66: frame_vm_group_bin_1396 (RW)
0x67: frame_vm_group_bin_17557 (RW)
0x68: frame_vm_group_bin_10412 (RW)
0x69: frame_vm_group_bin_3260 (RW)
0x6: frame_vm_group_bin_13719 (RW)
0x6a: frame_vm_group_bin_19330 (RW)
0x6b: frame_vm_group_bin_12156 (RW)
0x6c: frame_vm_group_bin_5058 (RW)
0x6d: frame_vm_group_bin_21155 (RW)
0x6e: frame_vm_group_bin_13978 (RW)
0x6f: frame_vm_group_bin_6796 (RW)
0x70: frame_vm_group_bin_22993 (RW)
0x71: frame_vm_group_bin_15810 (RW)
0x72: frame_vm_group_bin_8617 (RW)
0x73: frame_vm_group_bin_1429 (RW)
0x74: frame_vm_group_bin_17580 (RW)
0x75: frame_vm_group_bin_10440 (RW)
0x76: frame_vm_group_bin_3293 (RW)
0x77: frame_vm_group_bin_19363 (RW)
0x78: frame_vm_group_bin_14314 (RW)
0x79: frame_vm_group_bin_5092 (RW)
0x7: frame_vm_group_bin_6531 (RW)
0x7a: frame_vm_group_bin_21189 (RW)
0x7b: frame_vm_group_bin_14012 (RW)
0x7c: frame_vm_group_bin_6827 (RW)
0x7d: frame_vm_group_bin_23026 (RW)
0x7e: frame_vm_group_bin_15843 (RW)
0x7f: frame_vm_group_bin_8651 (RW)
0x80: frame_vm_group_bin_1463 (RW)
0x81: frame_vm_group_bin_17605 (RW)
0x82: frame_vm_group_bin_10474 (RW)
0x83: frame_vm_group_bin_3327 (RW)
0x84: frame_vm_group_bin_19397 (RW)
0x85: frame_vm_group_bin_12216 (RW)
0x86: frame_vm_group_bin_5126 (RW)
0x87: frame_vm_group_bin_21222 (RW)
0x88: frame_vm_group_bin_14045 (RW)
0x89: frame_vm_group_bin_13217 (RW)
0x8: frame_vm_group_bin_22728 (RW)
0x8a: frame_vm_group_bin_23059 (RW)
0x8b: frame_vm_group_bin_15876 (RW)
0x8c: frame_vm_group_bin_8685 (RW)
0x8d: frame_vm_group_bin_1496 (RW)
0x8e: frame_vm_group_bin_17636 (RW)
0x8f: frame_vm_group_bin_10507 (RW)
0x90: frame_vm_group_bin_3360 (RW)
0x91: frame_vm_group_bin_19429 (RW)
0x92: frame_vm_group_bin_12248 (RW)
0x93: frame_vm_group_bin_5159 (RW)
0x94: frame_vm_group_bin_21255 (RW)
0x95: frame_vm_group_bin_14078 (RW)
0x96: frame_vm_group_bin_6879 (RW)
0x97: frame_vm_group_bin_23092 (RW)
0x98: frame_vm_group_bin_15909 (RW)
0x99: frame_vm_group_bin_8718 (RW)
0x9: frame_vm_group_bin_15544 (RW)
0x9a: frame_vm_group_bin_1530 (RW)
0x9b: frame_vm_group_bin_17670 (RW)
0x9c: frame_vm_group_bin_10540 (RW)
0x9d: frame_vm_group_bin_3391 (RW)
0x9e: frame_vm_group_bin_19460 (RW)
0x9f: frame_vm_group_bin_12282 (RW)
0xa0: frame_vm_group_bin_5193 (RW)
0xa1: frame_vm_group_bin_21289 (RW)
0xa2: frame_vm_group_bin_14112 (RW)
0xa3: frame_vm_group_bin_22598 (RW)
0xa4: frame_vm_group_bin_23126 (RW)
0xa5: frame_vm_group_bin_15943 (RW)
0xa6: frame_vm_group_bin_8752 (RW)
0xa7: frame_vm_group_bin_1563 (RW)
0xa8: frame_vm_group_bin_17698 (RW)
0xa9: frame_vm_group_bin_10573 (RW)
0xa: frame_vm_group_bin_8354 (RW)
0xaa: frame_vm_group_bin_12512 (RW)
0xab: frame_vm_group_bin_19493 (RW)
0xac: frame_vm_group_bin_12315 (RW)
0xad: frame_vm_group_bin_5226 (RW)
0xae: frame_vm_group_bin_21321 (RW)
0xaf: frame_vm_group_bin_14145 (RW)
0xb0: frame_vm_group_bin_6933 (RW)
0xb1: frame_vm_group_bin_23158 (RW)
0xb2: frame_vm_group_bin_15976 (RW)
0xb3: frame_vm_group_bin_8785 (RW)
0xb4: frame_vm_group_bin_1596 (RW)
0xb5: frame_vm_group_bin_17723 (RW)
0xb6: frame_vm_group_bin_10606 (RW)
0xb7: frame_vm_group_bin_17259 (RW)
0xb8: frame_vm_group_bin_19526 (RW)
0xb9: frame_vm_group_bin_12347 (RW)
0xb: frame_vm_group_bin_1165 (RW)
0xba: frame_vm_group_bin_5260 (RW)
0xbb: frame_vm_group_bin_21354 (RW)
0xbc: frame_vm_group_bin_14179 (RW)
0xbd: frame_vm_group_bin_6966 (RW)
0xbe: frame_vm_group_bin_23191 (RW)
0xbf: frame_vm_group_bin_16012 (RW)
0xc0: frame_vm_group_bin_8819 (RW)
0xc1: frame_vm_group_bin_1630 (RW)
0xc2: frame_vm_group_bin_17751 (RW)
0xc3: frame_vm_group_bin_10640 (RW)
0xc4: frame_vm_group_bin_21895 (RW)
0xc5: frame_vm_group_bin_19560 (RW)
0xc6: frame_vm_group_bin_12381 (RW)
0xc7: frame_vm_group_bin_5293 (RW)
0xc8: frame_vm_group_bin_21387 (RW)
0xc9: frame_vm_group_bin_14211 (RW)
0xc: frame_vm_group_bin_17389 (RW)
0xca: frame_vm_group_bin_6998 (RW)
0xcb: frame_vm_group_bin_11821 (RW)
0xcc: frame_vm_group_bin_16045 (RW)
0xcd: frame_vm_group_bin_8852 (RW)
0xce: frame_vm_group_bin_1663 (RW)
0xcf: frame_vm_group_bin_17781 (RW)
0xd0: frame_vm_group_bin_10671 (RW)
0xd1: frame_vm_group_bin_3272 (RW)
0xd2: frame_vm_group_bin_19594 (RW)
0xd3: frame_vm_group_bin_12414 (RW)
0xd4: frame_vm_group_bin_5325 (RW)
0xd5: frame_vm_group_bin_21420 (RW)
0xd6: frame_vm_group_bin_14244 (RW)
0xd7: frame_vm_group_bin_7031 (RW)
0xd8: frame_vm_group_bin_23238 (RW)
0xd9: frame_vm_group_bin_16078 (RW)
0xd: frame_vm_group_bin_10187 (RW)
0xda: frame_vm_group_bin_8885 (RW)
0xdb: frame_vm_group_bin_1697 (RW)
0xdc: frame_vm_group_bin_17812 (RW)
0xdd: frame_vm_group_bin_10705 (RW)
0xde: frame_vm_group_bin_3520 (RW)
0xdf: frame_vm_group_bin_19628 (RW)
0xe0: frame_vm_group_bin_12447 (RW)
0xe1: frame_vm_group_bin_5357 (RW)
0xe2: frame_vm_group_bin_21453 (RW)
0xe3: frame_vm_group_bin_14277 (RW)
0xe4: frame_vm_group_bin_7063 (RW)
0xe5: frame_vm_group_bin_0008 (RW)
0xe6: frame_vm_group_bin_16111 (RW)
0xe7: frame_vm_group_bin_8917 (RW)
0xe8: frame_vm_group_bin_1729 (RW)
0xe9: frame_vm_group_bin_17841 (RW)
0xe: frame_vm_group_bin_3028 (RW)
0xea: frame_vm_group_bin_10737 (RW)
0xeb: frame_vm_group_bin_3551 (RW)
0xec: frame_vm_group_bin_5796 (RW)
0xed: frame_vm_group_bin_12479 (RW)
0xee: frame_vm_group_bin_5389 (RW)
0xef: frame_vm_group_bin_21485 (RW)
0xf0: frame_vm_group_bin_14308 (RW)
0xf1: frame_vm_group_bin_7095 (RW)
0xf2: frame_vm_group_bin_0026 (RW)
0xf3: frame_vm_group_bin_16142 (RW)
0xf4: frame_vm_group_bin_8949 (RW)
0xf5: frame_vm_group_bin_1761 (RW)
0xf6: frame_vm_group_bin_17867 (RW)
0xf7: frame_vm_group_bin_10770 (RW)
0xf8: frame_vm_group_bin_3583 (RW)
0xf9: frame_vm_group_bin_19684 (RW)
0xf: frame_vm_group_bin_19098 (RW)
0xfa: frame_vm_group_bin_12513 (RW)
0xfb: frame_vm_group_bin_5423 (RW)
0xfc: frame_vm_group_bin_21518 (RW)
0xfd: frame_vm_group_bin_14342 (RW)
0xfe: frame_vm_group_bin_7128 (RW)
0xff: frame_vm_group_bin_0049 (RW)
}
pt_vm_group_bin_0018 {
0x0: frame_vm_group_bin_12283 (RW)
0x100: frame_vm_group_bin_18291 (RW)
0x101: frame_vm_group_bin_11203 (RW)
0x102: frame_vm_group_bin_4018 (RW)
0x103: frame_vm_group_bin_20114 (RW)
0x104: frame_vm_group_bin_12915 (RW)
0x105: frame_vm_group_bin_5816 (RW)
0x106: frame_vm_group_bin_21951 (RW)
0x107: frame_vm_group_bin_14776 (RW)
0x108: frame_vm_group_bin_7560 (RW)
0x109: frame_vm_group_bin_0404 (RW)
0x10: frame_vm_group_bin_14146 (RW)
0x10a: frame_vm_group_bin_16591 (RW)
0x10b: frame_vm_group_bin_9380 (RW)
0x10c: frame_vm_group_bin_2225 (RW)
0x10d: frame_vm_group_bin_18324 (RW)
0x10e: frame_vm_group_bin_11236 (RW)
0x10f: frame_vm_group_bin_4051 (RW)
0x110: frame_vm_group_bin_20147 (RW)
0x111: frame_vm_group_bin_12947 (RW)
0x112: frame_vm_group_bin_5841 (RW)
0x113: frame_vm_group_bin_21984 (RW)
0x114: frame_vm_group_bin_14808 (RW)
0x115: frame_vm_group_bin_7593 (RW)
0x116: frame_vm_group_bin_0433 (RW)
0x117: frame_vm_group_bin_16623 (RW)
0x118: frame_vm_group_bin_9414 (RW)
0x119: frame_vm_group_bin_2254 (RW)
0x11: frame_vm_group_bin_6934 (RW)
0x11a: frame_vm_group_bin_18358 (RW)
0x11b: frame_vm_group_bin_11270 (RW)
0x11c: frame_vm_group_bin_4085 (RW)
0x11d: frame_vm_group_bin_20180 (RW)
0x11e: frame_vm_group_bin_12981 (RW)
0x11f: frame_vm_group_bin_5865 (RW)
0x120: frame_vm_group_bin_22017 (RW)
0x121: frame_vm_group_bin_14842 (RW)
0x122: frame_vm_group_bin_7627 (RW)
0x123: frame_vm_group_bin_0467 (RW)
0x124: frame_vm_group_bin_16657 (RW)
0x125: frame_vm_group_bin_9448 (RW)
0x126: frame_vm_group_bin_2288 (RW)
0x127: frame_vm_group_bin_18391 (RW)
0x128: frame_vm_group_bin_11303 (RW)
0x129: frame_vm_group_bin_4117 (RW)
0x12: frame_vm_group_bin_23159 (RW)
0x12a: frame_vm_group_bin_20212 (RW)
0x12b: frame_vm_group_bin_13016 (RW)
0x12c: frame_vm_group_bin_5891 (RW)
0x12d: frame_vm_group_bin_11196 (RW)
0x12e: frame_vm_group_bin_14875 (RW)
0x12f: frame_vm_group_bin_7660 (RW)
0x130: frame_vm_group_bin_0499 (RW)
0x131: frame_vm_group_bin_16690 (RW)
0x132: frame_vm_group_bin_9481 (RW)
0x133: frame_vm_group_bin_2321 (RW)
0x134: frame_vm_group_bin_18422 (RW)
0x135: frame_vm_group_bin_11336 (RW)
0x136: frame_vm_group_bin_4150 (RW)
0x137: frame_vm_group_bin_20245 (RW)
0x138: frame_vm_group_bin_13049 (RW)
0x139: frame_vm_group_bin_5917 (RW)
0x13: frame_vm_group_bin_15977 (RW)
0x13a: frame_vm_group_bin_22064 (RW)
0x13b: frame_vm_group_bin_14909 (RW)
0x13c: frame_vm_group_bin_7694 (RW)
0x13d: frame_vm_group_bin_0532 (RW)
0x13e: frame_vm_group_bin_16724 (RW)
0x13f: frame_vm_group_bin_9515 (RW)
0x140: frame_vm_group_bin_2355 (RW)
0x141: frame_vm_group_bin_18456 (RW)
0x142: frame_vm_group_bin_11368 (RW)
0x143: frame_vm_group_bin_4183 (RW)
0x144: frame_vm_group_bin_20278 (RW)
0x145: frame_vm_group_bin_13083 (RW)
0x146: frame_vm_group_bin_5941 (RW)
0x147: frame_vm_group_bin_22092 (RW)
0x148: frame_vm_group_bin_14942 (RW)
0x149: frame_vm_group_bin_7726 (RW)
0x14: frame_vm_group_bin_8786 (RW)
0x14a: frame_vm_group_bin_0563 (RW)
0x14b: frame_vm_group_bin_16757 (RW)
0x14c: frame_vm_group_bin_9548 (RW)
0x14d: frame_vm_group_bin_2388 (RW)
0x14e: frame_vm_group_bin_18483 (RW)
0x14f: frame_vm_group_bin_11400 (RW)
0x150: frame_vm_group_bin_4215 (RW)
0x151: frame_vm_group_bin_20311 (RW)
0x152: frame_vm_group_bin_13116 (RW)
0x153: frame_vm_group_bin_5966 (RW)
0x154: frame_vm_group_bin_22124 (RW)
0x155: frame_vm_group_bin_14975 (RW)
0x156: frame_vm_group_bin_7759 (RW)
0x157: frame_vm_group_bin_0595 (RW)
0x158: frame_vm_group_bin_16790 (RW)
0x159: frame_vm_group_bin_9581 (RW)
0x15: frame_vm_group_bin_1597 (RW)
0x15a: frame_vm_group_bin_2422 (RW)
0x15b: frame_vm_group_bin_18512 (RW)
0x15c: frame_vm_group_bin_11433 (RW)
0x15d: frame_vm_group_bin_4249 (RW)
0x15e: frame_vm_group_bin_20347 (RW)
0x15f: frame_vm_group_bin_13150 (RW)
0x160: frame_vm_group_bin_5995 (RW)
0x161: frame_vm_group_bin_22158 (RW)
0x162: frame_vm_group_bin_15009 (RW)
0x163: frame_vm_group_bin_7793 (RW)
0x164: frame_vm_group_bin_0627 (RW)
0x165: frame_vm_group_bin_16824 (RW)
0x166: frame_vm_group_bin_9615 (RW)
0x167: frame_vm_group_bin_2454 (RW)
0x168: frame_vm_group_bin_18537 (RW)
0x169: frame_vm_group_bin_11466 (RW)
0x16: frame_vm_group_bin_17724 (RW)
0x16a: frame_vm_group_bin_4282 (RW)
0x16b: frame_vm_group_bin_20380 (RW)
0x16c: frame_vm_group_bin_13183 (RW)
0x16d: frame_vm_group_bin_6026 (RW)
0x16e: frame_vm_group_bin_22191 (RW)
0x16f: frame_vm_group_bin_9747 (RW)
0x170: frame_vm_group_bin_7826 (RW)
0x171: frame_vm_group_bin_0661 (RW)
0x172: frame_vm_group_bin_16857 (RW)
0x173: frame_vm_group_bin_9648 (RW)
0x174: frame_vm_group_bin_2486 (RW)
0x175: frame_vm_group_bin_18563 (RW)
0x176: frame_vm_group_bin_11499 (RW)
0x177: frame_vm_group_bin_4315 (RW)
0x178: frame_vm_group_bin_20413 (RW)
0x179: frame_vm_group_bin_13216 (RW)
0x17: frame_vm_group_bin_10607 (RW)
0x17a: frame_vm_group_bin_6053 (RW)
0x17b: frame_vm_group_bin_22225 (RW)
0x17c: frame_vm_group_bin_15065 (RW)
0x17d: frame_vm_group_bin_7859 (RW)
0x17e: frame_vm_group_bin_0695 (RW)
0x17f: frame_vm_group_bin_10122 (RW)
0x180: frame_vm_group_bin_9681 (RW)
0x181: frame_vm_group_bin_2520 (RW)
0x182: frame_vm_group_bin_18597 (RW)
0x183: frame_vm_group_bin_11533 (RW)
0x184: frame_vm_group_bin_4351 (RW)
0x185: frame_vm_group_bin_20447 (RW)
0x186: frame_vm_group_bin_13250 (RW)
0x187: frame_vm_group_bin_6078 (RW)
0x188: frame_vm_group_bin_22258 (RW)
0x189: frame_vm_group_bin_15089 (RW)
0x18: frame_vm_group_bin_3438 (RW)
0x18a: frame_vm_group_bin_7892 (RW)
0x18b: frame_vm_group_bin_0728 (RW)
0x18c: frame_vm_group_bin_16922 (RW)
0x18d: frame_vm_group_bin_9714 (RW)
0x18e: frame_vm_group_bin_2553 (RW)
0x18f: frame_vm_group_bin_18630 (RW)
0x190: frame_vm_group_bin_9048 (RW)
0x191: frame_vm_group_bin_4384 (RW)
0x192: frame_vm_group_bin_20480 (RW)
0x193: frame_vm_group_bin_13283 (RW)
0x194: frame_vm_group_bin_6109 (RW)
0x195: frame_vm_group_bin_22290 (RW)
0x196: frame_vm_group_bin_15116 (RW)
0x197: frame_vm_group_bin_7925 (RW)
0x198: frame_vm_group_bin_0761 (RW)
0x199: frame_vm_group_bin_16955 (RW)
0x19: frame_vm_group_bin_19527 (RW)
0x19a: frame_vm_group_bin_9748 (RW)
0x19b: frame_vm_group_bin_2587 (RW)
0x19c: frame_vm_group_bin_18663 (RW)
0x19d: frame_vm_group_bin_11592 (RW)
0x19e: frame_vm_group_bin_4418 (RW)
0x19f: frame_vm_group_bin_20514 (RW)
0x1: frame_vm_group_bin_5194 (RW)
0x1a0: frame_vm_group_bin_13316 (RW)
0x1a1: frame_vm_group_bin_6141 (RW)
0x1a2: frame_vm_group_bin_22324 (RW)
0x1a3: frame_vm_group_bin_15140 (RW)
0x1a4: frame_vm_group_bin_7960 (RW)
0x1a5: frame_vm_group_bin_0795 (RW)
0x1a6: frame_vm_group_bin_16989 (RW)
0x1a7: frame_vm_group_bin_9781 (RW)
0x1a8: frame_vm_group_bin_2620 (RW)
0x1a9: frame_vm_group_bin_18696 (RW)
0x1a: frame_vm_group_bin_12349 (RW)
0x1aa: frame_vm_group_bin_11617 (RW)
0x1ab: frame_vm_group_bin_4451 (RW)
0x1ac: frame_vm_group_bin_20547 (RW)
0x1ad: frame_vm_group_bin_13349 (RW)
0x1ae: frame_vm_group_bin_6174 (RW)
0x1af: frame_vm_group_bin_22356 (RW)
0x1b0: frame_vm_group_bin_15172 (RW)
0x1b1: frame_vm_group_bin_7992 (RW)
0x1b2: frame_vm_group_bin_0827 (RW)
0x1b3: frame_vm_group_bin_17022 (RW)
0x1b4: frame_vm_group_bin_9814 (RW)
0x1b5: frame_vm_group_bin_2653 (RW)
0x1b6: frame_vm_group_bin_18728 (RW)
0x1b7: frame_vm_group_bin_11638 (RW)
0x1b8: frame_vm_group_bin_4484 (RW)
0x1b9: frame_vm_group_bin_20580 (RW)
0x1b: frame_vm_group_bin_5261 (RW)
0x1ba: frame_vm_group_bin_13381 (RW)
0x1bb: frame_vm_group_bin_17353 (RW)
0x1bc: frame_vm_group_bin_22390 (RW)
0x1bd: frame_vm_group_bin_15206 (RW)
0x1be: frame_vm_group_bin_8023 (RW)
0x1bf: frame_vm_group_bin_0861 (RW)
0x1c0: frame_vm_group_bin_17056 (RW)
0x1c1: frame_vm_group_bin_9848 (RW)
0x1c2: frame_vm_group_bin_2687 (RW)
0x1c3: frame_vm_group_bin_18760 (RW)
0x1c4: frame_vm_group_bin_11662 (RW)
0x1c5: frame_vm_group_bin_4518 (RW)
0x1c6: frame_vm_group_bin_20614 (RW)
0x1c7: frame_vm_group_bin_13414 (RW)
0x1c8: frame_vm_group_bin_6232 (RW)
0x1c9: frame_vm_group_bin_22422 (RW)
0x1c: frame_vm_group_bin_21355 (RW)
0x1ca: frame_vm_group_bin_15240 (RW)
0x1cb: frame_vm_group_bin_8051 (RW)
0x1cc: frame_vm_group_bin_0894 (RW)
0x1cd: frame_vm_group_bin_17089 (RW)
0x1ce: frame_vm_group_bin_9881 (RW)
0x1cf: frame_vm_group_bin_2720 (RW)
0x1d0: frame_vm_group_bin_18793 (RW)
0x1d1: frame_vm_group_bin_11686 (RW)
0x1d2: frame_vm_group_bin_4551 (RW)
0x1d3: frame_vm_group_bin_20647 (RW)
0x1d4: frame_vm_group_bin_13447 (RW)
0x1d5: frame_vm_group_bin_6263 (RW)
0x1d6: frame_vm_group_bin_22455 (RW)
0x1d7: frame_vm_group_bin_15273 (RW)
0x1d8: frame_vm_group_bin_22340 (RW)
0x1d9: frame_vm_group_bin_0927 (RW)
0x1d: frame_vm_group_bin_4996 (RW)
0x1da: frame_vm_group_bin_17123 (RW)
0x1db: frame_vm_group_bin_9914 (RW)
0x1dc: frame_vm_group_bin_2754 (RW)
0x1dd: frame_vm_group_bin_15155 (RW)
0x1de: frame_vm_group_bin_11715 (RW)
0x1df: frame_vm_group_bin_4580 (RW)
0x1e0: frame_vm_group_bin_20680 (RW)
0x1e1: frame_vm_group_bin_13481 (RW)
0x1e2: frame_vm_group_bin_6296 (RW)
0x1e3: frame_vm_group_bin_22489 (RW)
0x1e4: frame_vm_group_bin_15306 (RW)
0x1e5: frame_vm_group_bin_8115 (RW)
0x1e6: frame_vm_group_bin_0961 (RW)
0x1e7: frame_vm_group_bin_17155 (RW)
0x1e8: frame_vm_group_bin_9945 (RW)
0x1e9: frame_vm_group_bin_2787 (RW)
0x1e: frame_vm_group_bin_3538 (RW)
0x1ea: frame_vm_group_bin_18861 (RW)
0x1eb: frame_vm_group_bin_11739 (RW)
0x1ec: frame_vm_group_bin_4601 (RW)
0x1ed: frame_vm_group_bin_20713 (RW)
0x1ee: frame_vm_group_bin_13514 (RW)
0x1ef: frame_vm_group_bin_6328 (RW)
0x1f0: frame_vm_group_bin_22522 (RW)
0x1f1: frame_vm_group_bin_15339 (RW)
0x1f2: frame_vm_group_bin_8148 (RW)
0x1f3: frame_vm_group_bin_0994 (RW)
0x1f4: frame_vm_group_bin_17187 (RW)
0x1f5: frame_vm_group_bin_9978 (RW)
0x1f6: frame_vm_group_bin_2820 (RW)
0x1f7: frame_vm_group_bin_18894 (RW)
0x1f8: frame_vm_group_bin_11760 (RW)
0x1f9: frame_vm_group_bin_21634 (RW)
0x1f: frame_vm_group_bin_23192 (RW)
0x1fa: frame_vm_group_bin_20747 (RW)
0x1fb: frame_vm_group_bin_13548 (RW)
0x1fc: frame_vm_group_bin_6362 (RW)
0x1fd: frame_vm_group_bin_22555 (RW)
0x1fe: frame_vm_group_bin_15373 (RW)
0x1ff: frame_vm_group_bin_8182 (RW)
0x20: frame_vm_group_bin_16013 (RW)
0x21: frame_vm_group_bin_8820 (RW)
0x22: frame_vm_group_bin_1631 (RW)
0x23: frame_vm_group_bin_17752 (RW)
0x24: frame_vm_group_bin_10641 (RW)
0x25: frame_vm_group_bin_3464 (RW)
0x26: frame_vm_group_bin_19561 (RW)
0x27: frame_vm_group_bin_12382 (RW)
0x28: frame_vm_group_bin_5294 (RW)
0x29: frame_vm_group_bin_21388 (RW)
0x2: frame_vm_group_bin_21290 (RW)
0x2a: frame_vm_group_bin_14212 (RW)
0x2b: frame_vm_group_bin_6999 (RW)
0x2c: frame_vm_group_bin_6734 (RW)
0x2d: frame_vm_group_bin_16046 (RW)
0x2e: frame_vm_group_bin_8853 (RW)
0x2f: frame_vm_group_bin_1664 (RW)
0x30: frame_vm_group_bin_17782 (RW)
0x31: frame_vm_group_bin_10672 (RW)
0x32: frame_vm_group_bin_3490 (RW)
0x33: frame_vm_group_bin_19595 (RW)
0x34: frame_vm_group_bin_12415 (RW)
0x35: frame_vm_group_bin_5326 (RW)
0x36: frame_vm_group_bin_21421 (RW)
0x37: frame_vm_group_bin_14245 (RW)
0x38: frame_vm_group_bin_7032 (RW)
0x39: frame_vm_group_bin_11476 (RW)
0x3: frame_vm_group_bin_14113 (RW)
0x3a: frame_vm_group_bin_16080 (RW)
0x3b: frame_vm_group_bin_8886 (RW)
0x3c: frame_vm_group_bin_1698 (RW)
0x3d: frame_vm_group_bin_17813 (RW)
0x3e: frame_vm_group_bin_10706 (RW)
0x3f: frame_vm_group_bin_2847 (RW)
0x40: frame_vm_group_bin_19629 (RW)
0x41: frame_vm_group_bin_12448 (RW)
0x42: frame_vm_group_bin_5358 (RW)
0x43: frame_vm_group_bin_21454 (RW)
0x44: frame_vm_group_bin_14278 (RW)
0x45: frame_vm_group_bin_7064 (RW)
0x46: frame_vm_group_bin_0009 (RW)
0x47: frame_vm_group_bin_16112 (RW)
0x48: frame_vm_group_bin_8918 (RW)
0x49: frame_vm_group_bin_1730 (RW)
0x4: frame_vm_group_bin_6904 (RW)
0x4a: frame_vm_group_bin_17842 (RW)
0x4b: frame_vm_group_bin_10738 (RW)
0x4c: frame_vm_group_bin_3552 (RW)
0x4d: frame_vm_group_bin_6035 (RW)
0x4e: frame_vm_group_bin_12480 (RW)
0x4f: frame_vm_group_bin_5390 (RW)
0x50: frame_vm_group_bin_21486 (RW)
0x51: frame_vm_group_bin_14309 (RW)
0x52: frame_vm_group_bin_7096 (RW)
0x53: frame_vm_group_bin_0027 (RW)
0x54: frame_vm_group_bin_16143 (RW)
0x55: frame_vm_group_bin_8950 (RW)
0x56: frame_vm_group_bin_1762 (RW)
0x57: frame_vm_group_bin_17868 (RW)
0x58: frame_vm_group_bin_10771 (RW)
0x59: frame_vm_group_bin_3585 (RW)
0x5: frame_vm_group_bin_23127 (RW)
0x5a: frame_vm_group_bin_19686 (RW)
0x5b: frame_vm_group_bin_12514 (RW)
0x5c: frame_vm_group_bin_5424 (RW)
0x5d: frame_vm_group_bin_21519 (RW)
0x5e: frame_vm_group_bin_14343 (RW)
0x5f: frame_vm_group_bin_3561 (RW)
0x60: frame_vm_group_bin_0050 (RW)
0x61: frame_vm_group_bin_16177 (RW)
0x62: frame_vm_group_bin_8984 (RW)
0x63: frame_vm_group_bin_1796 (RW)
0x64: frame_vm_group_bin_17899 (RW)
0x65: frame_vm_group_bin_10804 (RW)
0x66: frame_vm_group_bin_3619 (RW)
0x67: frame_vm_group_bin_19719 (RW)
0x68: frame_vm_group_bin_12547 (RW)
0x69: frame_vm_group_bin_5456 (RW)
0x6: frame_vm_group_bin_15944 (RW)
0x6a: frame_vm_group_bin_21552 (RW)
0x6b: frame_vm_group_bin_14376 (RW)
0x6c: frame_vm_group_bin_7161 (RW)
0x6d: frame_vm_group_bin_0075 (RW)
0x6e: frame_vm_group_bin_5397 (RW)
0x6f: frame_vm_group_bin_9017 (RW)
0x70: frame_vm_group_bin_1829 (RW)
0x71: frame_vm_group_bin_17931 (RW)
0x72: frame_vm_group_bin_10837 (RW)
0x73: frame_vm_group_bin_3652 (RW)
0x74: frame_vm_group_bin_19752 (RW)
0x75: frame_vm_group_bin_12580 (RW)
0x76: frame_vm_group_bin_5488 (RW)
0x77: frame_vm_group_bin_21585 (RW)
0x78: frame_vm_group_bin_14409 (RW)
0x79: frame_vm_group_bin_7196 (RW)
0x7: frame_vm_group_bin_8753 (RW)
0x7a: frame_vm_group_bin_0102 (RW)
0x7b: frame_vm_group_bin_16236 (RW)
0x7c: frame_vm_group_bin_9051 (RW)
0x7d: frame_vm_group_bin_1863 (RW)
0x7e: frame_vm_group_bin_17963 (RW)
0x7f: frame_vm_group_bin_10870 (RW)
0x80: frame_vm_group_bin_3686 (RW)
0x81: frame_vm_group_bin_19786 (RW)
0x82: frame_vm_group_bin_12614 (RW)
0x83: frame_vm_group_bin_5521 (RW)
0x84: frame_vm_group_bin_21619 (RW)
0x85: frame_vm_group_bin_14443 (RW)
0x86: frame_vm_group_bin_7230 (RW)
0x87: frame_vm_group_bin_0126 (RW)
0x88: frame_vm_group_bin_16262 (RW)
0x89: frame_vm_group_bin_9084 (RW)
0x8: frame_vm_group_bin_1564 (RW)
0x8a: frame_vm_group_bin_1896 (RW)
0x8b: frame_vm_group_bin_17994 (RW)
0x8c: frame_vm_group_bin_10904 (RW)
0x8d: frame_vm_group_bin_3719 (RW)
0x8e: frame_vm_group_bin_19819 (RW)
0x8f: frame_vm_group_bin_12646 (RW)
0x90: frame_vm_group_bin_5554 (RW)
0x91: frame_vm_group_bin_21652 (RW)
0x92: frame_vm_group_bin_14476 (RW)
0x93: frame_vm_group_bin_7263 (RW)
0x94: frame_vm_group_bin_0147 (RW)
0x95: frame_vm_group_bin_16292 (RW)
0x96: frame_vm_group_bin_9117 (RW)
0x97: frame_vm_group_bin_1929 (RW)
0x98: frame_vm_group_bin_18027 (RW)
0x99: frame_vm_group_bin_10937 (RW)
0x9: frame_vm_group_bin_17699 (RW)
0x9a: frame_vm_group_bin_3753 (RW)
0x9b: frame_vm_group_bin_19853 (RW)
0x9c: frame_vm_group_bin_12673 (RW)
0x9d: frame_vm_group_bin_5587 (RW)
0x9e: frame_vm_group_bin_21685 (RW)
0x9f: frame_vm_group_bin_14511 (RW)
0xa0: frame_vm_group_bin_7296 (RW)
0xa1: frame_vm_group_bin_0171 (RW)
0xa2: frame_vm_group_bin_16325 (RW)
0xa3: frame_vm_group_bin_9150 (RW)
0xa4: frame_vm_group_bin_1962 (RW)
0xa5: frame_vm_group_bin_18060 (RW)
0xa6: frame_vm_group_bin_10970 (RW)
0xa7: frame_vm_group_bin_3785 (RW)
0xa8: frame_vm_group_bin_19885 (RW)
0xa9: frame_vm_group_bin_12696 (RW)
0xa: frame_vm_group_bin_10574 (RW)
0xaa: frame_vm_group_bin_5618 (RW)
0xab: frame_vm_group_bin_21718 (RW)
0xac: frame_vm_group_bin_14544 (RW)
0xad: frame_vm_group_bin_7329 (RW)
0xae: frame_vm_group_bin_0203 (RW)
0xaf: frame_vm_group_bin_16358 (RW)
0xb0: frame_vm_group_bin_9182 (RW)
0xb1: frame_vm_group_bin_1995 (RW)
0xb2: frame_vm_group_bin_18092 (RW)
0xb3: frame_vm_group_bin_11003 (RW)
0xb4: frame_vm_group_bin_3818 (RW)
0xb5: frame_vm_group_bin_19917 (RW)
0xb6: frame_vm_group_bin_12721 (RW)
0xb7: frame_vm_group_bin_5651 (RW)
0xb8: frame_vm_group_bin_21751 (RW)
0xb9: frame_vm_group_bin_14577 (RW)
0xb: frame_vm_group_bin_7431 (RW)
0xba: frame_vm_group_bin_7363 (RW)
0xbb: frame_vm_group_bin_0233 (RW)
0xbc: frame_vm_group_bin_16392 (RW)
0xbd: frame_vm_group_bin_9211 (RW)
0xbe: frame_vm_group_bin_2029 (RW)
0xbf: frame_vm_group_bin_18125 (RW)
0xc0: frame_vm_group_bin_11037 (RW)
0xc1: frame_vm_group_bin_3852 (RW)
0xc2: frame_vm_group_bin_19950 (RW)
0xc3: frame_vm_group_bin_12749 (RW)
0xc4: frame_vm_group_bin_5685 (RW)
0xc5: frame_vm_group_bin_21784 (RW)
0xc6: frame_vm_group_bin_14610 (RW)
0xc7: frame_vm_group_bin_7396 (RW)
0xc8: frame_vm_group_bin_0255 (RW)
0xc9: frame_vm_group_bin_16425 (RW)
0xc: frame_vm_group_bin_19494 (RW)
0xca: frame_vm_group_bin_9235 (RW)
0xcb: frame_vm_group_bin_2062 (RW)
0xcc: frame_vm_group_bin_18158 (RW)
0xcd: frame_vm_group_bin_11070 (RW)
0xce: frame_vm_group_bin_3885 (RW)
0xcf: frame_vm_group_bin_19983 (RW)
0xd0: frame_vm_group_bin_12782 (RW)
0xd1: frame_vm_group_bin_5718 (RW)
0xd2: frame_vm_group_bin_21818 (RW)
0xd3: frame_vm_group_bin_14643 (RW)
0xd4: frame_vm_group_bin_7429 (RW)
0xd5: frame_vm_group_bin_0279 (RW)
0xd6: frame_vm_group_bin_16458 (RW)
0xd7: frame_vm_group_bin_9258 (RW)
0xd8: frame_vm_group_bin_2095 (RW)
0xd9: frame_vm_group_bin_15079 (RW)
0xd: frame_vm_group_bin_12316 (RW)
0xda: frame_vm_group_bin_11104 (RW)
0xdb: frame_vm_group_bin_3919 (RW)
0xdc: frame_vm_group_bin_20015 (RW)
0xdd: frame_vm_group_bin_12816 (RW)
0xde: frame_vm_group_bin_5748 (RW)
0xdf: frame_vm_group_bin_21852 (RW)
0xe0: frame_vm_group_bin_14677 (RW)
0xe1: frame_vm_group_bin_7463 (RW)
0xe2: frame_vm_group_bin_0310 (RW)
0xe3: frame_vm_group_bin_16492 (RW)
0xe4: frame_vm_group_bin_9284 (RW)
0xe5: frame_vm_group_bin_2130 (RW)
0xe6: frame_vm_group_bin_18224 (RW)
0xe7: frame_vm_group_bin_11136 (RW)
0xe8: frame_vm_group_bin_3951 (RW)
0xe9: frame_vm_group_bin_20048 (RW)
0xe: frame_vm_group_bin_5227 (RW)
0xea: frame_vm_group_bin_12848 (RW)
0xeb: frame_vm_group_bin_5771 (RW)
0xec: frame_vm_group_bin_21885 (RW)
0xed: frame_vm_group_bin_14710 (RW)
0xee: frame_vm_group_bin_7496 (RW)
0xef: frame_vm_group_bin_0342 (RW)
0xf0: frame_vm_group_bin_16525 (RW)
0xf1: frame_vm_group_bin_9313 (RW)
0xf2: frame_vm_group_bin_2163 (RW)
0xf3: frame_vm_group_bin_18257 (RW)
0xf4: frame_vm_group_bin_11169 (RW)
0xf5: frame_vm_group_bin_3984 (RW)
0xf6: frame_vm_group_bin_20081 (RW)
0xf7: frame_vm_group_bin_12881 (RW)
0xf8: frame_vm_group_bin_5794 (RW)
0xf9: frame_vm_group_bin_21917 (RW)
0xf: frame_vm_group_bin_21322 (RW)
0xfa: frame_vm_group_bin_14743 (RW)
0xfb: frame_vm_group_bin_7529 (RW)
0xfc: frame_vm_group_bin_0374 (RW)
0xfd: frame_vm_group_bin_16558 (RW)
0xfe: frame_vm_group_bin_9347 (RW)
0xff: frame_vm_group_bin_2196 (RW)
}
pt_vm_group_bin_0020 {
0x0: frame_vm_group_bin_2495 (RW)
0x100: frame_vm_group_bin_8490 (RW)
0x101: frame_vm_group_bin_1298 (RW)
0x102: frame_vm_group_bin_17485 (RW)
0x103: frame_vm_group_bin_10323 (RW)
0x104: frame_vm_group_bin_3163 (RW)
0x105: frame_vm_group_bin_19232 (RW)
0x106: frame_vm_group_bin_12060 (RW)
0x107: frame_vm_group_bin_4961 (RW)
0x108: frame_vm_group_bin_21058 (RW)
0x109: frame_vm_group_bin_13880 (RW)
0x10: frame_vm_group_bin_4359 (RW)
0x10a: frame_vm_group_bin_6700 (RW)
0x10b: frame_vm_group_bin_22896 (RW)
0x10c: frame_vm_group_bin_15713 (RW)
0x10d: frame_vm_group_bin_8522 (RW)
0x10e: frame_vm_group_bin_1330 (RW)
0x10f: frame_vm_group_bin_17509 (RW)
0x110: frame_vm_group_bin_10356 (RW)
0x111: frame_vm_group_bin_3196 (RW)
0x112: frame_vm_group_bin_19265 (RW)
0x113: frame_vm_group_bin_12092 (RW)
0x114: frame_vm_group_bin_4993 (RW)
0x115: frame_vm_group_bin_21091 (RW)
0x116: frame_vm_group_bin_13913 (RW)
0x117: frame_vm_group_bin_6732 (RW)
0x118: frame_vm_group_bin_22929 (RW)
0x119: frame_vm_group_bin_15746 (RW)
0x11: frame_vm_group_bin_20455 (RW)
0x11a: frame_vm_group_bin_3459 (RW)
0x11b: frame_vm_group_bin_1366 (RW)
0x11c: frame_vm_group_bin_17538 (RW)
0x11d: frame_vm_group_bin_10389 (RW)
0x11e: frame_vm_group_bin_20999 (RW)
0x11f: frame_vm_group_bin_19299 (RW)
0x120: frame_vm_group_bin_12125 (RW)
0x121: frame_vm_group_bin_5027 (RW)
0x122: frame_vm_group_bin_21125 (RW)
0x123: frame_vm_group_bin_13947 (RW)
0x124: frame_vm_group_bin_6765 (RW)
0x125: frame_vm_group_bin_22962 (RW)
0x126: frame_vm_group_bin_15780 (RW)
0x127: frame_vm_group_bin_8587 (RW)
0x128: frame_vm_group_bin_1398 (RW)
0x129: frame_vm_group_bin_17559 (RW)
0x12: frame_vm_group_bin_13258 (RW)
0x12a: frame_vm_group_bin_10414 (RW)
0x12b: frame_vm_group_bin_3262 (RW)
0x12c: frame_vm_group_bin_19332 (RW)
0x12d: frame_vm_group_bin_12158 (RW)
0x12e: frame_vm_group_bin_5060 (RW)
0x12f: frame_vm_group_bin_21157 (RW)
0x130: frame_vm_group_bin_13980 (RW)
0x131: frame_vm_group_bin_6798 (RW)
0x132: frame_vm_group_bin_22995 (RW)
0x133: frame_vm_group_bin_15812 (RW)
0x134: frame_vm_group_bin_8619 (RW)
0x135: frame_vm_group_bin_1431 (RW)
0x136: frame_vm_group_bin_17582 (RW)
0x137: frame_vm_group_bin_10442 (RW)
0x138: frame_vm_group_bin_3295 (RW)
0x139: frame_vm_group_bin_19365 (RW)
0x13: frame_vm_group_bin_6086 (RW)
0x13a: frame_vm_group_bin_12188 (RW)
0x13b: frame_vm_group_bin_5095 (RW)
0x13c: frame_vm_group_bin_21191 (RW)
0x13d: frame_vm_group_bin_14014 (RW)
0x13e: frame_vm_group_bin_6829 (RW)
0x13f: frame_vm_group_bin_23028 (RW)
0x140: frame_vm_group_bin_15845 (RW)
0x141: frame_vm_group_bin_8653 (RW)
0x142: frame_vm_group_bin_1465 (RW)
0x143: frame_vm_group_bin_17607 (RW)
0x144: frame_vm_group_bin_10476 (RW)
0x145: frame_vm_group_bin_3329 (RW)
0x146: frame_vm_group_bin_19399 (RW)
0x147: frame_vm_group_bin_12218 (RW)
0x148: frame_vm_group_bin_5128 (RW)
0x149: frame_vm_group_bin_21224 (RW)
0x14: frame_vm_group_bin_22266 (RW)
0x14a: frame_vm_group_bin_14047 (RW)
0x14b: frame_vm_group_bin_6856 (RW)
0x14c: frame_vm_group_bin_23061 (RW)
0x14d: frame_vm_group_bin_15878 (RW)
0x14e: frame_vm_group_bin_8687 (RW)
0x14f: frame_vm_group_bin_1498 (RW)
0x150: frame_vm_group_bin_17638 (RW)
0x151: frame_vm_group_bin_10509 (RW)
0x152: frame_vm_group_bin_3362 (RW)
0x153: frame_vm_group_bin_19431 (RW)
0x154: frame_vm_group_bin_12250 (RW)
0x155: frame_vm_group_bin_5161 (RW)
0x156: frame_vm_group_bin_21257 (RW)
0x157: frame_vm_group_bin_14080 (RW)
0x158: frame_vm_group_bin_6881 (RW)
0x159: frame_vm_group_bin_23094 (RW)
0x15: frame_vm_group_bin_15094 (RW)
0x15a: frame_vm_group_bin_15912 (RW)
0x15b: frame_vm_group_bin_8721 (RW)
0x15c: frame_vm_group_bin_1532 (RW)
0x15d: frame_vm_group_bin_17672 (RW)
0x15e: frame_vm_group_bin_10542 (RW)
0x15f: frame_vm_group_bin_3393 (RW)
0x160: frame_vm_group_bin_19462 (RW)
0x161: frame_vm_group_bin_12284 (RW)
0x162: frame_vm_group_bin_5195 (RW)
0x163: frame_vm_group_bin_21291 (RW)
0x164: frame_vm_group_bin_14114 (RW)
0x165: frame_vm_group_bin_6905 (RW)
0x166: frame_vm_group_bin_23128 (RW)
0x167: frame_vm_group_bin_15945 (RW)
0x168: frame_vm_group_bin_8754 (RW)
0x169: frame_vm_group_bin_1565 (RW)
0x16: frame_vm_group_bin_7900 (RW)
0x16a: frame_vm_group_bin_17700 (RW)
0x16b: frame_vm_group_bin_10575 (RW)
0x16c: frame_vm_group_bin_3417 (RW)
0x16d: frame_vm_group_bin_19495 (RW)
0x16e: frame_vm_group_bin_12317 (RW)
0x16f: frame_vm_group_bin_5228 (RW)
0x170: frame_vm_group_bin_21323 (RW)
0x171: frame_vm_group_bin_14147 (RW)
0x172: frame_vm_group_bin_6935 (RW)
0x173: frame_vm_group_bin_23160 (RW)
0x174: frame_vm_group_bin_15978 (RW)
0x175: frame_vm_group_bin_8787 (RW)
0x176: frame_vm_group_bin_1598 (RW)
0x177: frame_vm_group_bin_17725 (RW)
0x178: frame_vm_group_bin_10608 (RW)
0x179: frame_vm_group_bin_3439 (RW)
0x17: frame_vm_group_bin_0736 (RW)
0x17a: frame_vm_group_bin_19529 (RW)
0x17b: frame_vm_group_bin_12350 (RW)
0x17c: frame_vm_group_bin_5262 (RW)
0x17d: frame_vm_group_bin_21356 (RW)
0x17e: frame_vm_group_bin_14180 (RW)
0x17f: frame_vm_group_bin_6967 (RW)
0x180: frame_vm_group_bin_23193 (RW)
0x181: frame_vm_group_bin_16014 (RW)
0x182: frame_vm_group_bin_8821 (RW)
0x183: frame_vm_group_bin_1632 (RW)
0x184: frame_vm_group_bin_17753 (RW)
0x185: frame_vm_group_bin_10642 (RW)
0x186: frame_vm_group_bin_3465 (RW)
0x187: frame_vm_group_bin_19562 (RW)
0x188: frame_vm_group_bin_12383 (RW)
0x189: frame_vm_group_bin_5295 (RW)
0x18: frame_vm_group_bin_16930 (RW)
0x18a: frame_vm_group_bin_21389 (RW)
0x18b: frame_vm_group_bin_14213 (RW)
0x18c: frame_vm_group_bin_7000 (RW)
0x18d: frame_vm_group_bin_1672 (RW)
0x18e: frame_vm_group_bin_16047 (RW)
0x18f: frame_vm_group_bin_8854 (RW)
0x190: frame_vm_group_bin_1665 (RW)
0x191: frame_vm_group_bin_17783 (RW)
0x192: frame_vm_group_bin_10673 (RW)
0x193: frame_vm_group_bin_3491 (RW)
0x194: frame_vm_group_bin_19596 (RW)
0x195: frame_vm_group_bin_12416 (RW)
0x196: frame_vm_group_bin_5327 (RW)
0x197: frame_vm_group_bin_21422 (RW)
0x198: frame_vm_group_bin_14246 (RW)
0x199: frame_vm_group_bin_7033 (RW)
0x19: frame_vm_group_bin_9722 (RW)
0x19a: frame_vm_group_bin_23240 (RW)
0x19b: frame_vm_group_bin_16081 (RW)
0x19c: frame_vm_group_bin_8887 (RW)
0x19d: frame_vm_group_bin_1699 (RW)
0x19e: frame_vm_group_bin_17814 (RW)
0x19f: frame_vm_group_bin_10707 (RW)
0x1: frame_vm_group_bin_18572 (RW)
0x1a0: frame_vm_group_bin_3521 (RW)
0x1a1: frame_vm_group_bin_19630 (RW)
0x1a2: frame_vm_group_bin_12449 (RW)
0x1a3: frame_vm_group_bin_5359 (RW)
0x1a4: frame_vm_group_bin_21455 (RW)
0x1a5: frame_vm_group_bin_14279 (RW)
0x1a6: frame_vm_group_bin_7065 (RW)
0x1a7: frame_vm_group_bin_0010 (RW)
0x1a8: frame_vm_group_bin_16113 (RW)
0x1a9: frame_vm_group_bin_8919 (RW)
0x1a: frame_vm_group_bin_2562 (RW)
0x1aa: frame_vm_group_bin_1731 (RW)
0x1ab: frame_vm_group_bin_17843 (RW)
0x1ac: frame_vm_group_bin_10739 (RW)
0x1ad: frame_vm_group_bin_3553 (RW)
0x1ae: frame_vm_group_bin_19658 (RW)
0x1af: frame_vm_group_bin_12481 (RW)
0x1b0: frame_vm_group_bin_5391 (RW)
0x1b1: frame_vm_group_bin_21487 (RW)
0x1b2: frame_vm_group_bin_14310 (RW)
0x1b3: frame_vm_group_bin_7097 (RW)
0x1b4: frame_vm_group_bin_0028 (RW)
0x1b5: frame_vm_group_bin_16144 (RW)
0x1b6: frame_vm_group_bin_8951 (RW)
0x1b7: frame_vm_group_bin_1763 (RW)
0x1b8: frame_vm_group_bin_17869 (RW)
0x1b9: frame_vm_group_bin_8508 (RW)
0x1b: frame_vm_group_bin_18638 (RW)
0x1ba: frame_vm_group_bin_3587 (RW)
0x1bb: frame_vm_group_bin_19687 (RW)
0x1bc: frame_vm_group_bin_12515 (RW)
0x1bd: frame_vm_group_bin_5425 (RW)
0x1be: frame_vm_group_bin_21520 (RW)
0x1bf: frame_vm_group_bin_14344 (RW)
0x1c0: frame_vm_group_bin_7129 (RW)
0x1c1: frame_vm_group_bin_0051 (RW)
0x1c2: frame_vm_group_bin_16178 (RW)
0x1c3: frame_vm_group_bin_8985 (RW)
0x1c4: frame_vm_group_bin_1797 (RW)
0x1c5: frame_vm_group_bin_17900 (RW)
0x1c6: frame_vm_group_bin_10805 (RW)
0x1c7: frame_vm_group_bin_3620 (RW)
0x1c8: frame_vm_group_bin_19720 (RW)
0x1c9: frame_vm_group_bin_12548 (RW)
0x1c: frame_vm_group_bin_11572 (RW)
0x1ca: frame_vm_group_bin_5457 (RW)
0x1cb: frame_vm_group_bin_21553 (RW)
0x1cc: frame_vm_group_bin_14377 (RW)
0x1cd: frame_vm_group_bin_7162 (RW)
0x1ce: frame_vm_group_bin_0076 (RW)
0x1cf: frame_vm_group_bin_16208 (RW)
0x1d0: frame_vm_group_bin_9018 (RW)
0x1d1: frame_vm_group_bin_1830 (RW)
0x1d2: frame_vm_group_bin_17932 (RW)
0x1d3: frame_vm_group_bin_10838 (RW)
0x1d4: frame_vm_group_bin_3653 (RW)
0x1d5: frame_vm_group_bin_19753 (RW)
0x1d6: frame_vm_group_bin_12581 (RW)
0x1d7: frame_vm_group_bin_5489 (RW)
0x1d8: frame_vm_group_bin_21586 (RW)
0x1d9: frame_vm_group_bin_14410 (RW)
0x1d: frame_vm_group_bin_4393 (RW)
0x1da: frame_vm_group_bin_7198 (RW)
0x1db: frame_vm_group_bin_0103 (RW)
0x1dc: frame_vm_group_bin_16237 (RW)
0x1dd: frame_vm_group_bin_9052 (RW)
0x1de: frame_vm_group_bin_1864 (RW)
0x1df: frame_vm_group_bin_17964 (RW)
0x1e0: frame_vm_group_bin_10871 (RW)
0x1e1: frame_vm_group_bin_3687 (RW)
0x1e2: frame_vm_group_bin_19787 (RW)
0x1e3: frame_vm_group_bin_12615 (RW)
0x1e4: frame_vm_group_bin_5522 (RW)
0x1e5: frame_vm_group_bin_21620 (RW)
0x1e6: frame_vm_group_bin_14444 (RW)
0x1e7: frame_vm_group_bin_7231 (RW)
0x1e8: frame_vm_group_bin_0127 (RW)
0x1e9: frame_vm_group_bin_16263 (RW)
0x1e: frame_vm_group_bin_20489 (RW)
0x1ea: frame_vm_group_bin_9085 (RW)
0x1eb: frame_vm_group_bin_1897 (RW)
0x1ec: frame_vm_group_bin_17995 (RW)
0x1ed: frame_vm_group_bin_10905 (RW)
0x1ee: frame_vm_group_bin_3720 (RW)
0x1ef: frame_vm_group_bin_19820 (RW)
0x1f0: frame_vm_group_bin_22906 (RW)
0x1f1: frame_vm_group_bin_5555 (RW)
0x1f2: frame_vm_group_bin_21653 (RW)
0x1f3: frame_vm_group_bin_14477 (RW)
0x1f4: frame_vm_group_bin_7264 (RW)
0x1f5: frame_vm_group_bin_0148 (RW)
0x1f6: frame_vm_group_bin_16293 (RW)
0x1f7: frame_vm_group_bin_9118 (RW)
0x1f8: frame_vm_group_bin_1930 (RW)
0x1f9: frame_vm_group_bin_18028 (RW)
0x1f: frame_vm_group_bin_13292 (RW)
0x1fa: frame_vm_group_bin_10939 (RW)
0x1fb: frame_vm_group_bin_3754 (RW)
0x1fc: frame_vm_group_bin_19854 (RW)
0x1fd: frame_vm_group_bin_12674 (RW)
0x1fe: frame_vm_group_bin_5588 (RW)
0x1ff: frame_vm_group_bin_21686 (RW)
0x20: frame_vm_group_bin_6117 (RW)
0x21: frame_vm_group_bin_22299 (RW)
0x22: frame_vm_group_bin_15124 (RW)
0x23: frame_vm_group_bin_7935 (RW)
0x24: frame_vm_group_bin_0770 (RW)
0x25: frame_vm_group_bin_16964 (RW)
0x26: frame_vm_group_bin_9756 (RW)
0x27: frame_vm_group_bin_2595 (RW)
0x28: frame_vm_group_bin_18671 (RW)
0x29: frame_vm_group_bin_11597 (RW)
0x2: frame_vm_group_bin_11508 (RW)
0x2a: frame_vm_group_bin_4426 (RW)
0x2b: frame_vm_group_bin_20522 (RW)
0x2c: frame_vm_group_bin_13324 (RW)
0x2d: frame_vm_group_bin_6149 (RW)
0x2e: frame_vm_group_bin_22332 (RW)
0x2f: frame_vm_group_bin_15147 (RW)
0x30: frame_vm_group_bin_7968 (RW)
0x31: frame_vm_group_bin_0803 (RW)
0x32: frame_vm_group_bin_16997 (RW)
0x33: frame_vm_group_bin_9789 (RW)
0x34: frame_vm_group_bin_2628 (RW)
0x35: frame_vm_group_bin_18703 (RW)
0x36: frame_vm_group_bin_11622 (RW)
0x37: frame_vm_group_bin_4459 (RW)
0x38: frame_vm_group_bin_20555 (RW)
0x39: frame_vm_group_bin_13357 (RW)
0x3: frame_vm_group_bin_4324 (RW)
0x3a: frame_vm_group_bin_6183 (RW)
0x3b: frame_vm_group_bin_22365 (RW)
0x3c: frame_vm_group_bin_15181 (RW)
0x3d: frame_vm_group_bin_8000 (RW)
0x3e: frame_vm_group_bin_0836 (RW)
0x3f: frame_vm_group_bin_17031 (RW)
0x40: frame_vm_group_bin_9823 (RW)
0x41: frame_vm_group_bin_2662 (RW)
0x42: frame_vm_group_bin_18735 (RW)
0x43: frame_vm_group_bin_11646 (RW)
0x44: frame_vm_group_bin_4493 (RW)
0x45: frame_vm_group_bin_20589 (RW)
0x46: frame_vm_group_bin_13389 (RW)
0x47: frame_vm_group_bin_6211 (RW)
0x48: frame_vm_group_bin_22398 (RW)
0x49: frame_vm_group_bin_15214 (RW)
0x4: frame_vm_group_bin_20422 (RW)
0x4a: frame_vm_group_bin_8028 (RW)
0x4b: frame_vm_group_bin_0869 (RW)
0x4c: frame_vm_group_bin_17064 (RW)
0x4d: frame_vm_group_bin_9856 (RW)
0x4e: frame_vm_group_bin_2695 (RW)
0x4f: frame_vm_group_bin_18768 (RW)
0x50: frame_vm_group_bin_11667 (RW)
0x51: frame_vm_group_bin_4526 (RW)
0x52: frame_vm_group_bin_20622 (RW)
0x53: frame_vm_group_bin_13422 (RW)
0x54: frame_vm_group_bin_6239 (RW)
0x55: frame_vm_group_bin_22430 (RW)
0x56: frame_vm_group_bin_15248 (RW)
0x57: frame_vm_group_bin_8058 (RW)
0x58: frame_vm_group_bin_0902 (RW)
0x59: frame_vm_group_bin_17097 (RW)
0x5: frame_vm_group_bin_13225 (RW)
0x5a: frame_vm_group_bin_9889 (RW)
0x5b: frame_vm_group_bin_2729 (RW)
0x5c: frame_vm_group_bin_18802 (RW)
0x5d: frame_vm_group_bin_11694 (RW)
0x5e: frame_vm_group_bin_4559 (RW)
0x5f: frame_vm_group_bin_20655 (RW)
0x60: frame_vm_group_bin_13456 (RW)
0x61: frame_vm_group_bin_6271 (RW)
0x62: frame_vm_group_bin_22464 (RW)
0x63: frame_vm_group_bin_15281 (RW)
0x64: frame_vm_group_bin_8091 (RW)
0x65: frame_vm_group_bin_0936 (RW)
0x66: frame_vm_group_bin_17131 (RW)
0x67: frame_vm_group_bin_9922 (RW)
0x68: frame_vm_group_bin_2762 (RW)
0x69: frame_vm_group_bin_18836 (RW)
0x6: frame_vm_group_bin_6060 (RW)
0x6a: frame_vm_group_bin_11722 (RW)
0x6b: frame_vm_group_bin_21307 (RW)
0x6c: frame_vm_group_bin_20688 (RW)
0x6d: frame_vm_group_bin_13489 (RW)
0x6e: frame_vm_group_bin_6304 (RW)
0x6f: frame_vm_group_bin_22497 (RW)
0x70: frame_vm_group_bin_15314 (RW)
0x71: frame_vm_group_bin_8123 (RW)
0x72: frame_vm_group_bin_0969 (RW)
0x73: frame_vm_group_bin_17163 (RW)
0x74: frame_vm_group_bin_9953 (RW)
0x75: frame_vm_group_bin_2795 (RW)
0x76: frame_vm_group_bin_18869 (RW)
0x77: frame_vm_group_bin_11744 (RW)
0x78: frame_vm_group_bin_4607 (RW)
0x79: frame_vm_group_bin_20721 (RW)
0x7: frame_vm_group_bin_22233 (RW)
0x7a: frame_vm_group_bin_13523 (RW)
0x7b: frame_vm_group_bin_6337 (RW)
0x7c: frame_vm_group_bin_22530 (RW)
0x7d: frame_vm_group_bin_15348 (RW)
0x7e: frame_vm_group_bin_8157 (RW)
0x7f: frame_vm_group_bin_1003 (RW)
0x80: frame_vm_group_bin_17194 (RW)
0x81: frame_vm_group_bin_9987 (RW)
0x82: frame_vm_group_bin_2829 (RW)
0x83: frame_vm_group_bin_18903 (RW)
0x84: frame_vm_group_bin_11768 (RW)
0x85: frame_vm_group_bin_4634 (RW)
0x86: frame_vm_group_bin_20755 (RW)
0x87: frame_vm_group_bin_13556 (RW)
0x88: frame_vm_group_bin_6370 (RW)
0x89: frame_vm_group_bin_22563 (RW)
0x8: frame_vm_group_bin_15070 (RW)
0x8a: frame_vm_group_bin_15381 (RW)
0x8b: frame_vm_group_bin_8190 (RW)
0x8c: frame_vm_group_bin_20604 (RW)
0x8d: frame_vm_group_bin_17227 (RW)
0x8e: frame_vm_group_bin_10020 (RW)
0x8f: frame_vm_group_bin_2861 (RW)
0x90: frame_vm_group_bin_18936 (RW)
0x91: frame_vm_group_bin_11793 (RW)
0x92: frame_vm_group_bin_4667 (RW)
0x93: frame_vm_group_bin_20788 (RW)
0x94: frame_vm_group_bin_13589 (RW)
0x95: frame_vm_group_bin_6400 (RW)
0x96: frame_vm_group_bin_22596 (RW)
0x97: frame_vm_group_bin_15414 (RW)
0x98: frame_vm_group_bin_8223 (RW)
0x99: frame_vm_group_bin_1050 (RW)
0x9: frame_vm_group_bin_7867 (RW)
0x9a: frame_vm_group_bin_17260 (RW)
0x9b: frame_vm_group_bin_10054 (RW)
0x9c: frame_vm_group_bin_2897 (RW)
0x9d: frame_vm_group_bin_18968 (RW)
0x9e: frame_vm_group_bin_11826 (RW)
0x9f: frame_vm_group_bin_4699 (RW)
0xa0: frame_vm_group_bin_20821 (RW)
0xa1: frame_vm_group_bin_13623 (RW)
0xa2: frame_vm_group_bin_6433 (RW)
0xa3: frame_vm_group_bin_22630 (RW)
0xa4: frame_vm_group_bin_15448 (RW)
0xa5: frame_vm_group_bin_8257 (RW)
0xa6: frame_vm_group_bin_1074 (RW)
0xa7: frame_vm_group_bin_17293 (RW)
0xa8: frame_vm_group_bin_10087 (RW)
0xa9: frame_vm_group_bin_2930 (RW)
0xa: frame_vm_group_bin_0703 (RW)
0xaa: frame_vm_group_bin_19000 (RW)
0xab: frame_vm_group_bin_11856 (RW)
0xac: frame_vm_group_bin_4731 (RW)
0xad: frame_vm_group_bin_19874 (RW)
0xae: frame_vm_group_bin_13655 (RW)
0xaf: frame_vm_group_bin_6466 (RW)
0xb0: frame_vm_group_bin_22663 (RW)
0xb1: frame_vm_group_bin_15481 (RW)
0xb2: frame_vm_group_bin_8289 (RW)
0xb3: frame_vm_group_bin_1101 (RW)
0xb4: frame_vm_group_bin_17326 (RW)
0xb5: frame_vm_group_bin_10120 (RW)
0xb6: frame_vm_group_bin_2963 (RW)
0xb7: frame_vm_group_bin_19033 (RW)
0xb8: frame_vm_group_bin_11884 (RW)
0xb9: frame_vm_group_bin_4764 (RW)
0xb: frame_vm_group_bin_16897 (RW)
0xba: frame_vm_group_bin_20876 (RW)
0xbb: frame_vm_group_bin_13689 (RW)
0xbc: frame_vm_group_bin_6500 (RW)
0xbd: frame_vm_group_bin_22697 (RW)
0xbe: frame_vm_group_bin_15514 (RW)
0xbf: frame_vm_group_bin_8323 (RW)
0xc0: frame_vm_group_bin_1134 (RW)
0xc1: frame_vm_group_bin_17359 (RW)
0xc2: frame_vm_group_bin_10156 (RW)
0xc3: frame_vm_group_bin_2997 (RW)
0xc4: frame_vm_group_bin_19067 (RW)
0xc5: frame_vm_group_bin_11908 (RW)
0xc6: frame_vm_group_bin_4798 (RW)
0xc7: frame_vm_group_bin_20903 (RW)
0xc8: frame_vm_group_bin_13721 (RW)
0xc9: frame_vm_group_bin_6533 (RW)
0xc: frame_vm_group_bin_9689 (RW)
0xca: frame_vm_group_bin_22730 (RW)
0xcb: frame_vm_group_bin_15546 (RW)
0xcc: frame_vm_group_bin_8356 (RW)
0xcd: frame_vm_group_bin_1167 (RW)
0xce: frame_vm_group_bin_19151 (RW)
0xcf: frame_vm_group_bin_10189 (RW)
0xd0: frame_vm_group_bin_3030 (RW)
0xd1: frame_vm_group_bin_19100 (RW)
0xd2: frame_vm_group_bin_11938 (RW)
0xd3: frame_vm_group_bin_4830 (RW)
0xd4: frame_vm_group_bin_20931 (RW)
0xd5: frame_vm_group_bin_13754 (RW)
0xd6: frame_vm_group_bin_6566 (RW)
0xd7: frame_vm_group_bin_22762 (RW)
0xd8: frame_vm_group_bin_15579 (RW)
0xd9: frame_vm_group_bin_8389 (RW)
0xd: frame_vm_group_bin_2528 (RW)
0xda: frame_vm_group_bin_1201 (RW)
0xdb: frame_vm_group_bin_0528 (RW)
0xdc: frame_vm_group_bin_10223 (RW)
0xdd: frame_vm_group_bin_3064 (RW)
0xde: frame_vm_group_bin_19132 (RW)
0xdf: frame_vm_group_bin_11969 (RW)
0xe0: frame_vm_group_bin_4864 (RW)
0xe1: frame_vm_group_bin_20959 (RW)
0xe2: frame_vm_group_bin_13789 (RW)
0xe3: frame_vm_group_bin_6600 (RW)
0xe4: frame_vm_group_bin_22796 (RW)
0xe5: frame_vm_group_bin_15613 (RW)
0xe6: frame_vm_group_bin_8423 (RW)
0xe7: frame_vm_group_bin_1234 (RW)
0xe8: frame_vm_group_bin_17442 (RW)
0xe9: frame_vm_group_bin_10256 (RW)
0xe: frame_vm_group_bin_18605 (RW)
0xea: frame_vm_group_bin_3097 (RW)
0xeb: frame_vm_group_bin_19165 (RW)
0xec: frame_vm_group_bin_12001 (RW)
0xed: frame_vm_group_bin_4897 (RW)
0xee: frame_vm_group_bin_20990 (RW)
0xef: frame_vm_group_bin_18449 (RW)
0xf0: frame_vm_group_bin_6633 (RW)
0xf1: frame_vm_group_bin_22829 (RW)
0xf2: frame_vm_group_bin_15646 (RW)
0xf3: frame_vm_group_bin_8456 (RW)
0xf4: frame_vm_group_bin_1266 (RW)
0xf5: frame_vm_group_bin_17464 (RW)
0xf6: frame_vm_group_bin_10289 (RW)
0xf7: frame_vm_group_bin_3129 (RW)
0xf8: frame_vm_group_bin_19198 (RW)
0xf9: frame_vm_group_bin_12031 (RW)
0xf: frame_vm_group_bin_11541 (RW)
0xfa: frame_vm_group_bin_2727 (RW)
0xfb: frame_vm_group_bin_21024 (RW)
0xfc: frame_vm_group_bin_13851 (RW)
0xfd: frame_vm_group_bin_6667 (RW)
0xfe: frame_vm_group_bin_22863 (RW)
0xff: frame_vm_group_bin_15680 (RW)
}
pt_vm_group_bin_0022 {
0x0: frame_vm_group_bin_21428 (RW)
0x100: frame_vm_group_bin_4156 (RW)
0x101: frame_vm_group_bin_20252 (RW)
0x102: frame_vm_group_bin_13056 (RW)
0x103: frame_vm_group_bin_5923 (RW)
0x104: frame_vm_group_bin_11690 (RW)
0x105: frame_vm_group_bin_14915 (RW)
0x106: frame_vm_group_bin_7700 (RW)
0x107: frame_vm_group_bin_0538 (RW)
0x108: frame_vm_group_bin_16730 (RW)
0x109: frame_vm_group_bin_9521 (RW)
0x10: frame_vm_group_bin_0011 (RW)
0x10a: frame_vm_group_bin_2361 (RW)
0x10b: frame_vm_group_bin_18461 (RW)
0x10c: frame_vm_group_bin_11374 (RW)
0x10d: frame_vm_group_bin_4189 (RW)
0x10e: frame_vm_group_bin_20284 (RW)
0x10f: frame_vm_group_bin_13089 (RW)
0x110: frame_vm_group_bin_5945 (RW)
0x111: frame_vm_group_bin_22097 (RW)
0x112: frame_vm_group_bin_14948 (RW)
0x113: frame_vm_group_bin_7732 (RW)
0x114: frame_vm_group_bin_0569 (RW)
0x115: frame_vm_group_bin_16763 (RW)
0x116: frame_vm_group_bin_9554 (RW)
0x117: frame_vm_group_bin_2394 (RW)
0x118: frame_vm_group_bin_18488 (RW)
0x119: frame_vm_group_bin_11406 (RW)
0x11: frame_vm_group_bin_16118 (RW)
0x11a: frame_vm_group_bin_4222 (RW)
0x11b: frame_vm_group_bin_20320 (RW)
0x11c: frame_vm_group_bin_13123 (RW)
0x11d: frame_vm_group_bin_5970 (RW)
0x11e: frame_vm_group_bin_22131 (RW)
0x11f: frame_vm_group_bin_14982 (RW)
0x120: frame_vm_group_bin_7766 (RW)
0x121: frame_vm_group_bin_0602 (RW)
0x122: frame_vm_group_bin_16797 (RW)
0x123: frame_vm_group_bin_9588 (RW)
0x124: frame_vm_group_bin_2427 (RW)
0x125: frame_vm_group_bin_11006 (RW)
0x126: frame_vm_group_bin_11439 (RW)
0x127: frame_vm_group_bin_4255 (RW)
0x128: frame_vm_group_bin_20353 (RW)
0x129: frame_vm_group_bin_13156 (RW)
0x12: frame_vm_group_bin_8924 (RW)
0x12a: frame_vm_group_bin_6001 (RW)
0x12b: frame_vm_group_bin_22164 (RW)
0x12c: frame_vm_group_bin_15015 (RW)
0x12d: frame_vm_group_bin_7799 (RW)
0x12e: frame_vm_group_bin_0633 (RW)
0x12f: frame_vm_group_bin_16830 (RW)
0x130: frame_vm_group_bin_9621 (RW)
0x131: frame_vm_group_bin_2460 (RW)
0x132: frame_vm_group_bin_15651 (RW)
0x133: frame_vm_group_bin_11472 (RW)
0x134: frame_vm_group_bin_4288 (RW)
0x135: frame_vm_group_bin_20386 (RW)
0x136: frame_vm_group_bin_13189 (RW)
0x137: frame_vm_group_bin_6032 (RW)
0x138: frame_vm_group_bin_22197 (RW)
0x139: frame_vm_group_bin_15043 (RW)
0x13: frame_vm_group_bin_1736 (RW)
0x13a: frame_vm_group_bin_7832 (RW)
0x13b: frame_vm_group_bin_0668 (RW)
0x13c: frame_vm_group_bin_16864 (RW)
0x13d: frame_vm_group_bin_9655 (RW)
0x13e: frame_vm_group_bin_2493 (RW)
0x13f: frame_vm_group_bin_18570 (RW)
0x140: frame_vm_group_bin_11506 (RW)
0x141: frame_vm_group_bin_4322 (RW)
0x142: frame_vm_group_bin_20420 (RW)
0x143: frame_vm_group_bin_13223 (RW)
0x144: frame_vm_group_bin_6058 (RW)
0x145: frame_vm_group_bin_22231 (RW)
0x146: frame_vm_group_bin_10291 (RW)
0x147: frame_vm_group_bin_7865 (RW)
0x148: frame_vm_group_bin_0701 (RW)
0x149: frame_vm_group_bin_16895 (RW)
0x14: frame_vm_group_bin_17847 (RW)
0x14a: frame_vm_group_bin_9687 (RW)
0x14b: frame_vm_group_bin_2526 (RW)
0x14c: frame_vm_group_bin_18603 (RW)
0x14d: frame_vm_group_bin_11539 (RW)
0x14e: frame_vm_group_bin_4357 (RW)
0x14f: frame_vm_group_bin_20453 (RW)
0x150: frame_vm_group_bin_13256 (RW)
0x151: frame_vm_group_bin_6084 (RW)
0x152: frame_vm_group_bin_22264 (RW)
0x153: frame_vm_group_bin_14953 (RW)
0x154: frame_vm_group_bin_7898 (RW)
0x155: frame_vm_group_bin_0734 (RW)
0x156: frame_vm_group_bin_16928 (RW)
0x157: frame_vm_group_bin_9720 (RW)
0x158: frame_vm_group_bin_2559 (RW)
0x159: frame_vm_group_bin_18636 (RW)
0x15: frame_vm_group_bin_10744 (RW)
0x15a: frame_vm_group_bin_11570 (RW)
0x15b: frame_vm_group_bin_4391 (RW)
0x15c: frame_vm_group_bin_20487 (RW)
0x15d: frame_vm_group_bin_13290 (RW)
0x15e: frame_vm_group_bin_6115 (RW)
0x15f: frame_vm_group_bin_22297 (RW)
0x160: frame_vm_group_bin_19576 (RW)
0x161: frame_vm_group_bin_7933 (RW)
0x162: frame_vm_group_bin_0768 (RW)
0x163: frame_vm_group_bin_16962 (RW)
0x164: frame_vm_group_bin_9754 (RW)
0x165: frame_vm_group_bin_2593 (RW)
0x166: frame_vm_group_bin_18669 (RW)
0x167: frame_vm_group_bin_9558 (RW)
0x168: frame_vm_group_bin_4424 (RW)
0x169: frame_vm_group_bin_20520 (RW)
0x16: frame_vm_group_bin_3558 (RW)
0x16a: frame_vm_group_bin_13322 (RW)
0x16b: frame_vm_group_bin_6147 (RW)
0x16c: frame_vm_group_bin_22330 (RW)
0x16d: frame_vm_group_bin_15145 (RW)
0x16e: frame_vm_group_bin_7966 (RW)
0x16f: frame_vm_group_bin_0801 (RW)
0x170: frame_vm_group_bin_16995 (RW)
0x171: frame_vm_group_bin_9787 (RW)
0x172: frame_vm_group_bin_2626 (RW)
0x173: frame_vm_group_bin_15674 (RW)
0x174: frame_vm_group_bin_14223 (RW)
0x175: frame_vm_group_bin_4457 (RW)
0x176: frame_vm_group_bin_20553 (RW)
0x177: frame_vm_group_bin_13355 (RW)
0x178: frame_vm_group_bin_6180 (RW)
0x179: frame_vm_group_bin_22362 (RW)
0x17: frame_vm_group_bin_16717 (RW)
0x17a: frame_vm_group_bin_15179 (RW)
0x17b: frame_vm_group_bin_7998 (RW)
0x17c: frame_vm_group_bin_0834 (RW)
0x17d: frame_vm_group_bin_17029 (RW)
0x17e: frame_vm_group_bin_9821 (RW)
0x17f: frame_vm_group_bin_2660 (RW)
0x180: frame_vm_group_bin_18733 (RW)
0x181: frame_vm_group_bin_11644 (RW)
0x182: frame_vm_group_bin_4491 (RW)
0x183: frame_vm_group_bin_20587 (RW)
0x184: frame_vm_group_bin_13387 (RW)
0x185: frame_vm_group_bin_6209 (RW)
0x186: frame_vm_group_bin_22396 (RW)
0x187: frame_vm_group_bin_15212 (RW)
0x188: frame_vm_group_bin_8861 (RW)
0x189: frame_vm_group_bin_0867 (RW)
0x18: frame_vm_group_bin_12486 (RW)
0x18a: frame_vm_group_bin_17062 (RW)
0x18b: frame_vm_group_bin_9854 (RW)
0x18c: frame_vm_group_bin_2693 (RW)
0x18d: frame_vm_group_bin_18766 (RW)
0x18e: frame_vm_group_bin_11665 (RW)
0x18f: frame_vm_group_bin_4524 (RW)
0x190: frame_vm_group_bin_20620 (RW)
0x191: frame_vm_group_bin_13420 (RW)
0x192: frame_vm_group_bin_6237 (RW)
0x193: frame_vm_group_bin_22428 (RW)
0x194: frame_vm_group_bin_15246 (RW)
0x195: frame_vm_group_bin_8056 (RW)
0x196: frame_vm_group_bin_0900 (RW)
0x197: frame_vm_group_bin_17095 (RW)
0x198: frame_vm_group_bin_9887 (RW)
0x199: frame_vm_group_bin_2726 (RW)
0x19: frame_vm_group_bin_5396 (RW)
0x19a: frame_vm_group_bin_18800 (RW)
0x19b: frame_vm_group_bin_11692 (RW)
0x19c: frame_vm_group_bin_4557 (RW)
0x19d: frame_vm_group_bin_20653 (RW)
0x19e: frame_vm_group_bin_13454 (RW)
0x19f: frame_vm_group_bin_6269 (RW)
0x1: frame_vm_group_bin_14252 (RW)
0x1a0: frame_vm_group_bin_22462 (RW)
0x1a1: frame_vm_group_bin_15279 (RW)
0x1a2: frame_vm_group_bin_8089 (RW)
0x1a3: frame_vm_group_bin_0934 (RW)
0x1a4: frame_vm_group_bin_17129 (RW)
0x1a5: frame_vm_group_bin_9920 (RW)
0x1a6: frame_vm_group_bin_2760 (RW)
0x1a7: frame_vm_group_bin_18834 (RW)
0x1a8: frame_vm_group_bin_11720 (RW)
0x1a9: frame_vm_group_bin_8129 (RW)
0x1a: frame_vm_group_bin_21493 (RW)
0x1aa: frame_vm_group_bin_20686 (RW)
0x1ab: frame_vm_group_bin_13487 (RW)
0x1ac: frame_vm_group_bin_6302 (RW)
0x1ad: frame_vm_group_bin_22495 (RW)
0x1ae: frame_vm_group_bin_15312 (RW)
0x1af: frame_vm_group_bin_8121 (RW)
0x1b0: frame_vm_group_bin_0967 (RW)
0x1b1: frame_vm_group_bin_17161 (RW)
0x1b2: frame_vm_group_bin_9951 (RW)
0x1b3: frame_vm_group_bin_2793 (RW)
0x1b4: frame_vm_group_bin_18867 (RW)
0x1b5: frame_vm_group_bin_11742 (RW)
0x1b6: frame_vm_group_bin_4605 (RW)
0x1b7: frame_vm_group_bin_20719 (RW)
0x1b8: frame_vm_group_bin_13520 (RW)
0x1b9: frame_vm_group_bin_6334 (RW)
0x1b: frame_vm_group_bin_14316 (RW)
0x1ba: frame_vm_group_bin_22528 (RW)
0x1bb: frame_vm_group_bin_15346 (RW)
0x1bc: frame_vm_group_bin_8155 (RW)
0x1bd: frame_vm_group_bin_1001 (RW)
0x1be: frame_vm_group_bin_17192 (RW)
0x1bf: frame_vm_group_bin_9985 (RW)
0x1c0: frame_vm_group_bin_2827 (RW)
0x1c1: frame_vm_group_bin_18901 (RW)
0x1c2: frame_vm_group_bin_11766 (RW)
0x1c3: frame_vm_group_bin_4632 (RW)
0x1c4: frame_vm_group_bin_20753 (RW)
0x1c5: frame_vm_group_bin_13554 (RW)
0x1c6: frame_vm_group_bin_6368 (RW)
0x1c7: frame_vm_group_bin_22561 (RW)
0x1c8: frame_vm_group_bin_15379 (RW)
0x1c9: frame_vm_group_bin_8188 (RW)
0x1c: frame_vm_group_bin_7103 (RW)
0x1ca: frame_vm_group_bin_7408 (RW)
0x1cb: frame_vm_group_bin_17225 (RW)
0x1cc: frame_vm_group_bin_10018 (RW)
0x1cd: frame_vm_group_bin_2859 (RW)
0x1ce: frame_vm_group_bin_18934 (RW)
0x1cf: frame_vm_group_bin_11791 (RW)
0x1d0: frame_vm_group_bin_4665 (RW)
0x1d1: frame_vm_group_bin_20786 (RW)
0x1d2: frame_vm_group_bin_13587 (RW)
0x1d3: frame_vm_group_bin_6398 (RW)
0x1d4: frame_vm_group_bin_22594 (RW)
0x1d5: frame_vm_group_bin_15412 (RW)
0x1d6: frame_vm_group_bin_8221 (RW)
0x1d7: frame_vm_group_bin_12073 (RW)
0x1d8: frame_vm_group_bin_17257 (RW)
0x1d9: frame_vm_group_bin_10051 (RW)
0x1d: frame_vm_group_bin_0031 (RW)
0x1da: frame_vm_group_bin_2895 (RW)
0x1db: frame_vm_group_bin_18966 (RW)
0x1dc: frame_vm_group_bin_11824 (RW)
0x1dd: frame_vm_group_bin_3515 (RW)
0x1de: frame_vm_group_bin_2072 (RW)
0x1df: frame_vm_group_bin_13621 (RW)
0x1e0: frame_vm_group_bin_6431 (RW)
0x1e1: frame_vm_group_bin_22628 (RW)
0x1e2: frame_vm_group_bin_15446 (RW)
0x1e3: frame_vm_group_bin_8255 (RW)
0x1e4: frame_vm_group_bin_16815 (RW)
0x1e5: frame_vm_group_bin_17291 (RW)
0x1e6: frame_vm_group_bin_10085 (RW)
0x1e7: frame_vm_group_bin_2928 (RW)
0x1e8: frame_vm_group_bin_18998 (RW)
0x1e9: frame_vm_group_bin_11854 (RW)
0x1e: frame_vm_group_bin_16150 (RW)
0x1ea: frame_vm_group_bin_4729 (RW)
0x1eb: frame_vm_group_bin_20850 (RW)
0x1ec: frame_vm_group_bin_13653 (RW)
0x1ed: frame_vm_group_bin_6464 (RW)
0x1ee: frame_vm_group_bin_22661 (RW)
0x1ef: frame_vm_group_bin_15479 (RW)
0x1f0: frame_vm_group_bin_8287 (RW)
0x1f1: frame_vm_group_bin_1099 (RW)
0x1f2: frame_vm_group_bin_17324 (RW)
0x1f3: frame_vm_group_bin_10118 (RW)
0x1f4: frame_vm_group_bin_2961 (RW)
0x1f5: frame_vm_group_bin_19031 (RW)
0x1f6: frame_vm_group_bin_11882 (RW)
0x1f7: frame_vm_group_bin_4762 (RW)
0x1f8: frame_vm_group_bin_20873 (RW)
0x1f9: frame_vm_group_bin_13686 (RW)
0x1f: frame_vm_group_bin_8957 (RW)
0x1fa: frame_vm_group_bin_6498 (RW)
0x1fb: frame_vm_group_bin_22695 (RW)
0x1fc: frame_vm_group_bin_15512 (RW)
0x1fd: frame_vm_group_bin_8321 (RW)
0x1fe: frame_vm_group_bin_1132 (RW)
0x1ff: frame_vm_group_bin_1339 (RW)
0x20: frame_vm_group_bin_1769 (RW)
0x21: frame_vm_group_bin_17874 (RW)
0x22: frame_vm_group_bin_10777 (RW)
0x23: frame_vm_group_bin_3592 (RW)
0x24: frame_vm_group_bin_19692 (RW)
0x25: frame_vm_group_bin_12520 (RW)
0x26: frame_vm_group_bin_5430 (RW)
0x27: frame_vm_group_bin_21525 (RW)
0x28: frame_vm_group_bin_14349 (RW)
0x29: frame_vm_group_bin_7134 (RW)
0x2: frame_vm_group_bin_7039 (RW)
0x2a: frame_vm_group_bin_0054 (RW)
0x2b: frame_vm_group_bin_16183 (RW)
0x2c: frame_vm_group_bin_8990 (RW)
0x2d: frame_vm_group_bin_1802 (RW)
0x2e: frame_vm_group_bin_17905 (RW)
0x2f: frame_vm_group_bin_10810 (RW)
0x30: frame_vm_group_bin_3625 (RW)
0x31: frame_vm_group_bin_19725 (RW)
0x32: frame_vm_group_bin_12553 (RW)
0x33: frame_vm_group_bin_5462 (RW)
0x34: frame_vm_group_bin_21558 (RW)
0x35: frame_vm_group_bin_14382 (RW)
0x36: frame_vm_group_bin_7167 (RW)
0x37: frame_vm_group_bin_0080 (RW)
0x38: frame_vm_group_bin_16213 (RW)
0x39: frame_vm_group_bin_9023 (RW)
0x3: frame_vm_group_bin_7243 (RW)
0x3a: frame_vm_group_bin_1836 (RW)
0x3b: frame_vm_group_bin_17937 (RW)
0x3c: frame_vm_group_bin_10844 (RW)
0x3d: frame_vm_group_bin_3659 (RW)
0x3e: frame_vm_group_bin_19759 (RW)
0x3f: frame_vm_group_bin_12587 (RW)
0x40: frame_vm_group_bin_5495 (RW)
0x41: frame_vm_group_bin_21592 (RW)
0x42: frame_vm_group_bin_14416 (RW)
0x43: frame_vm_group_bin_7203 (RW)
0x44: frame_vm_group_bin_0106 (RW)
0x45: frame_vm_group_bin_5881 (RW)
0x46: frame_vm_group_bin_9057 (RW)
0x47: frame_vm_group_bin_1869 (RW)
0x48: frame_vm_group_bin_17969 (RW)
0x49: frame_vm_group_bin_10876 (RW)
0x4: frame_vm_group_bin_16086 (RW)
0x4a: frame_vm_group_bin_3692 (RW)
0x4b: frame_vm_group_bin_19792 (RW)
0x4c: frame_vm_group_bin_12620 (RW)
0x4d: frame_vm_group_bin_5527 (RW)
0x4e: frame_vm_group_bin_21625 (RW)
0x4f: frame_vm_group_bin_14449 (RW)
0x50: frame_vm_group_bin_7236 (RW)
0x51: frame_vm_group_bin_0129 (RW)
0x52: frame_vm_group_bin_16267 (RW)
0x53: frame_vm_group_bin_9090 (RW)
0x54: frame_vm_group_bin_1902 (RW)
0x55: frame_vm_group_bin_18000 (RW)
0x56: frame_vm_group_bin_10910 (RW)
0x57: frame_vm_group_bin_3725 (RW)
0x58: frame_vm_group_bin_19825 (RW)
0x59: frame_vm_group_bin_12651 (RW)
0x5: frame_vm_group_bin_8892 (RW)
0x5a: frame_vm_group_bin_5561 (RW)
0x5b: frame_vm_group_bin_21659 (RW)
0x5c: frame_vm_group_bin_14483 (RW)
0x5d: frame_vm_group_bin_7270 (RW)
0x5e: frame_vm_group_bin_0151 (RW)
0x5f: frame_vm_group_bin_16299 (RW)
0x60: frame_vm_group_bin_9124 (RW)
0x61: frame_vm_group_bin_1936 (RW)
0x62: frame_vm_group_bin_18034 (RW)
0x63: frame_vm_group_bin_10944 (RW)
0x64: frame_vm_group_bin_3759 (RW)
0x65: frame_vm_group_bin_19859 (RW)
0x66: frame_vm_group_bin_5213 (RW)
0x67: frame_vm_group_bin_5593 (RW)
0x68: frame_vm_group_bin_21691 (RW)
0x69: frame_vm_group_bin_14517 (RW)
0x6: frame_vm_group_bin_1704 (RW)
0x6a: frame_vm_group_bin_7302 (RW)
0x6b: frame_vm_group_bin_0177 (RW)
0x6c: frame_vm_group_bin_16331 (RW)
0x6d: frame_vm_group_bin_9156 (RW)
0x6e: frame_vm_group_bin_1968 (RW)
0x6f: frame_vm_group_bin_18066 (RW)
0x70: frame_vm_group_bin_10976 (RW)
0x71: frame_vm_group_bin_3791 (RW)
0x72: frame_vm_group_bin_19891 (RW)
0x73: frame_vm_group_bin_9841 (RW)
0x74: frame_vm_group_bin_5624 (RW)
0x75: frame_vm_group_bin_21724 (RW)
0x76: frame_vm_group_bin_14550 (RW)
0x77: frame_vm_group_bin_7335 (RW)
0x78: frame_vm_group_bin_0209 (RW)
0x79: frame_vm_group_bin_16364 (RW)
0x7: frame_vm_group_bin_17819 (RW)
0x7a: frame_vm_group_bin_9188 (RW)
0x7b: frame_vm_group_bin_2002 (RW)
0x7c: frame_vm_group_bin_20222 (RW)
0x7d: frame_vm_group_bin_11010 (RW)
0x7e: frame_vm_group_bin_3825 (RW)
0x7f: frame_vm_group_bin_15958 (RW)
0x80: frame_vm_group_bin_14505 (RW)
0x81: frame_vm_group_bin_5658 (RW)
0x82: frame_vm_group_bin_21758 (RW)
0x83: frame_vm_group_bin_14584 (RW)
0x84: frame_vm_group_bin_7369 (RW)
0x85: frame_vm_group_bin_0237 (RW)
0x86: frame_vm_group_bin_16398 (RW)
0x87: frame_vm_group_bin_4509 (RW)
0x88: frame_vm_group_bin_2035 (RW)
0x89: frame_vm_group_bin_18131 (RW)
0x8: frame_vm_group_bin_10712 (RW)
0x8a: frame_vm_group_bin_11043 (RW)
0x8b: frame_vm_group_bin_3858 (RW)
0x8c: frame_vm_group_bin_19956 (RW)
0x8d: frame_vm_group_bin_12755 (RW)
0x8e: frame_vm_group_bin_5691 (RW)
0x8f: frame_vm_group_bin_21790 (RW)
0x90: frame_vm_group_bin_14616 (RW)
0x91: frame_vm_group_bin_7402 (RW)
0x92: frame_vm_group_bin_0258 (RW)
0x93: frame_vm_group_bin_16431 (RW)
0x94: frame_vm_group_bin_9144 (RW)
0x95: frame_vm_group_bin_2068 (RW)
0x96: frame_vm_group_bin_18164 (RW)
0x97: frame_vm_group_bin_11076 (RW)
0x98: frame_vm_group_bin_3891 (RW)
0x99: frame_vm_group_bin_1955 (RW)
0x9: frame_vm_group_bin_3526 (RW)
0x9a: frame_vm_group_bin_12789 (RW)
0x9b: frame_vm_group_bin_5725 (RW)
0x9c: frame_vm_group_bin_21825 (RW)
0x9d: frame_vm_group_bin_14650 (RW)
0x9e: frame_vm_group_bin_7436 (RW)
0x9f: frame_vm_group_bin_0285 (RW)
0xa0: frame_vm_group_bin_16465 (RW)
0xa1: frame_vm_group_bin_13782 (RW)
0xa2: frame_vm_group_bin_2102 (RW)
0xa3: frame_vm_group_bin_18197 (RW)
0xa4: frame_vm_group_bin_11110 (RW)
0xa5: frame_vm_group_bin_3925 (RW)
0xa6: frame_vm_group_bin_20021 (RW)
0xa7: frame_vm_group_bin_12821 (RW)
0xa8: frame_vm_group_bin_3775 (RW)
0xa9: frame_vm_group_bin_21858 (RW)
0xa: frame_vm_group_bin_19635 (RW)
0xaa: frame_vm_group_bin_14683 (RW)
0xab: frame_vm_group_bin_7469 (RW)
0xac: frame_vm_group_bin_0316 (RW)
0xad: frame_vm_group_bin_16498 (RW)
0xae: frame_vm_group_bin_18424 (RW)
0xaf: frame_vm_group_bin_2136 (RW)
0xb0: frame_vm_group_bin_18230 (RW)
0xb1: frame_vm_group_bin_11142 (RW)
0xb2: frame_vm_group_bin_3957 (RW)
0xb3: frame_vm_group_bin_20054 (RW)
0xb4: frame_vm_group_bin_12854 (RW)
0xb5: frame_vm_group_bin_8414 (RW)
0xb6: frame_vm_group_bin_21891 (RW)
0xb7: frame_vm_group_bin_14716 (RW)
0xb8: frame_vm_group_bin_7502 (RW)
0xb9: frame_vm_group_bin_0347 (RW)
0xb: frame_vm_group_bin_12454 (RW)
0xba: frame_vm_group_bin_16532 (RW)
0xbb: frame_vm_group_bin_9320 (RW)
0xbc: frame_vm_group_bin_2170 (RW)
0xbd: frame_vm_group_bin_18264 (RW)
0xbe: frame_vm_group_bin_11176 (RW)
0xbf: frame_vm_group_bin_3991 (RW)
0xc0: frame_vm_group_bin_20088 (RW)
0xc1: frame_vm_group_bin_12888 (RW)
0xc2: frame_vm_group_bin_13051 (RW)
0xc3: frame_vm_group_bin_21924 (RW)
0xc4: frame_vm_group_bin_14749 (RW)
0xc5: frame_vm_group_bin_7534 (RW)
0xc6: frame_vm_group_bin_0380 (RW)
0xc7: frame_vm_group_bin_16564 (RW)
0xc8: frame_vm_group_bin_9353 (RW)
0xc9: frame_vm_group_bin_2202 (RW)
0xc: frame_vm_group_bin_5364 (RW)
0xca: frame_vm_group_bin_18297 (RW)
0xcb: frame_vm_group_bin_11209 (RW)
0xcc: frame_vm_group_bin_4024 (RW)
0xcd: frame_vm_group_bin_20120 (RW)
0xce: frame_vm_group_bin_12921 (RW)
0xcf: frame_vm_group_bin_5819 (RW)
0xd0: frame_vm_group_bin_21957 (RW)
0xd1: frame_vm_group_bin_14781 (RW)
0xd2: frame_vm_group_bin_7566 (RW)
0xd3: frame_vm_group_bin_0408 (RW)
0xd4: frame_vm_group_bin_10610 (RW)
0xd5: frame_vm_group_bin_9386 (RW)
0xd6: frame_vm_group_bin_2229 (RW)
0xd7: frame_vm_group_bin_18330 (RW)
0xd8: frame_vm_group_bin_11242 (RW)
0xd9: frame_vm_group_bin_4057 (RW)
0xd: frame_vm_group_bin_21460 (RW)
0xda: frame_vm_group_bin_20154 (RW)
0xdb: frame_vm_group_bin_12954 (RW)
0xdc: frame_vm_group_bin_5845 (RW)
0xdd: frame_vm_group_bin_21991 (RW)
0xde: frame_vm_group_bin_14815 (RW)
0xdf: frame_vm_group_bin_7600 (RW)
0xe0: frame_vm_group_bin_0440 (RW)
0xe1: frame_vm_group_bin_16630 (RW)
0xe2: frame_vm_group_bin_9421 (RW)
0xe3: frame_vm_group_bin_2261 (RW)
0xe4: frame_vm_group_bin_18364 (RW)
0xe5: frame_vm_group_bin_11276 (RW)
0xe6: frame_vm_group_bin_4091 (RW)
0xe7: frame_vm_group_bin_20185 (RW)
0xe8: frame_vm_group_bin_12987 (RW)
0xe9: frame_vm_group_bin_5870 (RW)
0xe: frame_vm_group_bin_14284 (RW)
0xea: frame_vm_group_bin_22022 (RW)
0xeb: frame_vm_group_bin_14848 (RW)
0xec: frame_vm_group_bin_7633 (RW)
0xed: frame_vm_group_bin_0473 (RW)
0xee: frame_vm_group_bin_16663 (RW)
0xef: frame_vm_group_bin_9454 (RW)
0xf0: frame_vm_group_bin_2294 (RW)
0xf1: frame_vm_group_bin_18396 (RW)
0xf2: frame_vm_group_bin_11309 (RW)
0xf3: frame_vm_group_bin_4123 (RW)
0xf4: frame_vm_group_bin_20218 (RW)
0xf5: frame_vm_group_bin_13022 (RW)
0xf6: frame_vm_group_bin_5895 (RW)
0xf7: frame_vm_group_bin_6962 (RW)
0xf8: frame_vm_group_bin_14881 (RW)
0xf9: frame_vm_group_bin_7666 (RW)
0xf: frame_vm_group_bin_7070 (RW)
0xfa: frame_vm_group_bin_0506 (RW)
0xfb: frame_vm_group_bin_1247 (RW)
0xfc: frame_vm_group_bin_9488 (RW)
0xfd: frame_vm_group_bin_2328 (RW)
0xfe: frame_vm_group_bin_18429 (RW)
0xff: frame_vm_group_bin_18799 (RW)
}
pt_vm_group_bin_0024 {
0x0: frame_vm_group_bin_13764 (RW)
0x100: frame_vm_group_bin_19761 (RW)
0x101: frame_vm_group_bin_12589 (RW)
0x102: frame_vm_group_bin_5497 (RW)
0x103: frame_vm_group_bin_21594 (RW)
0x104: frame_vm_group_bin_14418 (RW)
0x105: frame_vm_group_bin_7205 (RW)
0x106: frame_vm_group_bin_0108 (RW)
0x107: frame_vm_group_bin_16242 (RW)
0x108: frame_vm_group_bin_9059 (RW)
0x109: frame_vm_group_bin_1871 (RW)
0x10: frame_vm_group_bin_15621 (RW)
0x10a: frame_vm_group_bin_17971 (RW)
0x10b: frame_vm_group_bin_10878 (RW)
0x10c: frame_vm_group_bin_3694 (RW)
0x10d: frame_vm_group_bin_19794 (RW)
0x10e: frame_vm_group_bin_12622 (RW)
0x10f: frame_vm_group_bin_5529 (RW)
0x110: frame_vm_group_bin_21627 (RW)
0x111: frame_vm_group_bin_14451 (RW)
0x112: frame_vm_group_bin_7238 (RW)
0x113: frame_vm_group_bin_1812 (RW)
0x114: frame_vm_group_bin_16269 (RW)
0x115: frame_vm_group_bin_9092 (RW)
0x116: frame_vm_group_bin_1904 (RW)
0x117: frame_vm_group_bin_18002 (RW)
0x118: frame_vm_group_bin_10912 (RW)
0x119: frame_vm_group_bin_3727 (RW)
0x11: frame_vm_group_bin_8431 (RW)
0x11a: frame_vm_group_bin_19828 (RW)
0x11b: frame_vm_group_bin_12654 (RW)
0x11c: frame_vm_group_bin_5563 (RW)
0x11d: frame_vm_group_bin_21661 (RW)
0x11e: frame_vm_group_bin_14485 (RW)
0x11f: frame_vm_group_bin_7272 (RW)
0x120: frame_vm_group_bin_0153 (RW)
0x121: frame_vm_group_bin_16301 (RW)
0x122: frame_vm_group_bin_9126 (RW)
0x123: frame_vm_group_bin_1938 (RW)
0x124: frame_vm_group_bin_18036 (RW)
0x125: frame_vm_group_bin_10946 (RW)
0x126: frame_vm_group_bin_3761 (RW)
0x127: frame_vm_group_bin_19861 (RW)
0x128: frame_vm_group_bin_12678 (RW)
0x129: frame_vm_group_bin_5595 (RW)
0x12: frame_vm_group_bin_1242 (RW)
0x12a: frame_vm_group_bin_21693 (RW)
0x12b: frame_vm_group_bin_14519 (RW)
0x12c: frame_vm_group_bin_7304 (RW)
0x12d: frame_vm_group_bin_0179 (RW)
0x12e: frame_vm_group_bin_16333 (RW)
0x12f: frame_vm_group_bin_9158 (RW)
0x130: frame_vm_group_bin_1970 (RW)
0x131: frame_vm_group_bin_18068 (RW)
0x132: frame_vm_group_bin_10978 (RW)
0x133: frame_vm_group_bin_3793 (RW)
0x134: frame_vm_group_bin_19893 (RW)
0x135: frame_vm_group_bin_12702 (RW)
0x136: frame_vm_group_bin_5626 (RW)
0x137: frame_vm_group_bin_21726 (RW)
0x138: frame_vm_group_bin_14552 (RW)
0x139: frame_vm_group_bin_7337 (RW)
0x13: frame_vm_group_bin_17448 (RW)
0x13a: frame_vm_group_bin_0212 (RW)
0x13b: frame_vm_group_bin_16367 (RW)
0x13c: frame_vm_group_bin_9190 (RW)
0x13d: frame_vm_group_bin_2004 (RW)
0x13e: frame_vm_group_bin_10099 (RW)
0x13f: frame_vm_group_bin_11012 (RW)
0x140: frame_vm_group_bin_3827 (RW)
0x141: frame_vm_group_bin_19925 (RW)
0x142: frame_vm_group_bin_12729 (RW)
0x143: frame_vm_group_bin_5660 (RW)
0x144: frame_vm_group_bin_21760 (RW)
0x145: frame_vm_group_bin_14586 (RW)
0x146: frame_vm_group_bin_7371 (RW)
0x147: frame_vm_group_bin_0239 (RW)
0x148: frame_vm_group_bin_16400 (RW)
0x149: frame_vm_group_bin_9217 (RW)
0x14: frame_vm_group_bin_10264 (RW)
0x14a: frame_vm_group_bin_2037 (RW)
0x14b: frame_vm_group_bin_18133 (RW)
0x14c: frame_vm_group_bin_11045 (RW)
0x14d: frame_vm_group_bin_3860 (RW)
0x14e: frame_vm_group_bin_19958 (RW)
0x14f: frame_vm_group_bin_12757 (RW)
0x150: frame_vm_group_bin_5693 (RW)
0x151: frame_vm_group_bin_21792 (RW)
0x152: frame_vm_group_bin_14618 (RW)
0x153: frame_vm_group_bin_7404 (RW)
0x154: frame_vm_group_bin_0260 (RW)
0x155: frame_vm_group_bin_16433 (RW)
0x156: frame_vm_group_bin_9241 (RW)
0x157: frame_vm_group_bin_2070 (RW)
0x158: frame_vm_group_bin_18166 (RW)
0x159: frame_vm_group_bin_11078 (RW)
0x15: frame_vm_group_bin_3105 (RW)
0x15a: frame_vm_group_bin_3894 (RW)
0x15b: frame_vm_group_bin_15118 (RW)
0x15c: frame_vm_group_bin_12791 (RW)
0x15d: frame_vm_group_bin_5727 (RW)
0x15e: frame_vm_group_bin_21827 (RW)
0x15f: frame_vm_group_bin_14652 (RW)
0x160: frame_vm_group_bin_7438 (RW)
0x161: frame_vm_group_bin_0287 (RW)
0x162: frame_vm_group_bin_16467 (RW)
0x163: frame_vm_group_bin_9265 (RW)
0x164: frame_vm_group_bin_2104 (RW)
0x165: frame_vm_group_bin_18199 (RW)
0x166: frame_vm_group_bin_11112 (RW)
0x167: frame_vm_group_bin_3927 (RW)
0x168: frame_vm_group_bin_20023 (RW)
0x169: frame_vm_group_bin_12823 (RW)
0x16: frame_vm_group_bin_19173 (RW)
0x16a: frame_vm_group_bin_16956 (RW)
0x16b: frame_vm_group_bin_21860 (RW)
0x16c: frame_vm_group_bin_14685 (RW)
0x16d: frame_vm_group_bin_7471 (RW)
0x16e: frame_vm_group_bin_0318 (RW)
0x16f: frame_vm_group_bin_16500 (RW)
0x170: frame_vm_group_bin_9291 (RW)
0x171: frame_vm_group_bin_2138 (RW)
0x172: frame_vm_group_bin_18232 (RW)
0x173: frame_vm_group_bin_11144 (RW)
0x174: frame_vm_group_bin_3959 (RW)
0x175: frame_vm_group_bin_20056 (RW)
0x176: frame_vm_group_bin_12856 (RW)
0x177: frame_vm_group_bin_5777 (RW)
0x178: frame_vm_group_bin_21893 (RW)
0x179: frame_vm_group_bin_14718 (RW)
0x17: frame_vm_group_bin_12009 (RW)
0x17a: frame_vm_group_bin_17329 (RW)
0x17b: frame_vm_group_bin_0350 (RW)
0x17c: frame_vm_group_bin_16534 (RW)
0x17d: frame_vm_group_bin_9322 (RW)
0x17e: frame_vm_group_bin_2172 (RW)
0x17f: frame_vm_group_bin_18266 (RW)
0x180: frame_vm_group_bin_11178 (RW)
0x181: frame_vm_group_bin_3993 (RW)
0x182: frame_vm_group_bin_20090 (RW)
0x183: frame_vm_group_bin_12890 (RW)
0x184: frame_vm_group_bin_5800 (RW)
0x185: frame_vm_group_bin_21926 (RW)
0x186: frame_vm_group_bin_14751 (RW)
0x187: frame_vm_group_bin_7536 (RW)
0x188: frame_vm_group_bin_0382 (RW)
0x189: frame_vm_group_bin_16566 (RW)
0x18: frame_vm_group_bin_4905 (RW)
0x18a: frame_vm_group_bin_9355 (RW)
0x18b: frame_vm_group_bin_2203 (RW)
0x18c: frame_vm_group_bin_18299 (RW)
0x18d: frame_vm_group_bin_11211 (RW)
0x18e: frame_vm_group_bin_4026 (RW)
0x18f: frame_vm_group_bin_20122 (RW)
0x190: frame_vm_group_bin_12923 (RW)
0x191: frame_vm_group_bin_5821 (RW)
0x192: frame_vm_group_bin_21959 (RW)
0x193: frame_vm_group_bin_14783 (RW)
0x194: frame_vm_group_bin_7568 (RW)
0x195: frame_vm_group_bin_0410 (RW)
0x196: frame_vm_group_bin_16598 (RW)
0x197: frame_vm_group_bin_9388 (RW)
0x198: frame_vm_group_bin_2231 (RW)
0x199: frame_vm_group_bin_18332 (RW)
0x19: frame_vm_group_bin_20998 (RW)
0x19a: frame_vm_group_bin_11245 (RW)
0x19b: frame_vm_group_bin_4060 (RW)
0x19c: frame_vm_group_bin_15136 (RW)
0x19d: frame_vm_group_bin_12956 (RW)
0x19e: frame_vm_group_bin_5847 (RW)
0x19f: frame_vm_group_bin_21993 (RW)
0x1: frame_vm_group_bin_6575 (RW)
0x1a0: frame_vm_group_bin_14817 (RW)
0x1a1: frame_vm_group_bin_7602 (RW)
0x1a2: frame_vm_group_bin_0442 (RW)
0x1a3: frame_vm_group_bin_16632 (RW)
0x1a4: frame_vm_group_bin_9423 (RW)
0x1a5: frame_vm_group_bin_2263 (RW)
0x1a6: frame_vm_group_bin_18366 (RW)
0x1a7: frame_vm_group_bin_11278 (RW)
0x1a8: frame_vm_group_bin_4093 (RW)
0x1a9: frame_vm_group_bin_20187 (RW)
0x1a: frame_vm_group_bin_13829 (RW)
0x1aa: frame_vm_group_bin_12989 (RW)
0x1ab: frame_vm_group_bin_5872 (RW)
0x1ac: frame_vm_group_bin_15510 (RW)
0x1ad: frame_vm_group_bin_14850 (RW)
0x1ae: frame_vm_group_bin_7635 (RW)
0x1af: frame_vm_group_bin_0475 (RW)
0x1b0: frame_vm_group_bin_16665 (RW)
0x1b1: frame_vm_group_bin_9456 (RW)
0x1b2: frame_vm_group_bin_2296 (RW)
0x1b3: frame_vm_group_bin_18398 (RW)
0x1b4: frame_vm_group_bin_11311 (RW)
0x1b5: frame_vm_group_bin_4125 (RW)
0x1b6: frame_vm_group_bin_20220 (RW)
0x1b7: frame_vm_group_bin_13024 (RW)
0x1b8: frame_vm_group_bin_5897 (RW)
0x1b9: frame_vm_group_bin_20153 (RW)
0x1b: frame_vm_group_bin_6642 (RW)
0x1ba: frame_vm_group_bin_14884 (RW)
0x1bb: frame_vm_group_bin_7669 (RW)
0x1bc: frame_vm_group_bin_0508 (RW)
0x1bd: frame_vm_group_bin_16698 (RW)
0x1be: frame_vm_group_bin_9490 (RW)
0x1bf: frame_vm_group_bin_2330 (RW)
0x1c0: frame_vm_group_bin_18431 (RW)
0x1c1: frame_vm_group_bin_11343 (RW)
0x1c2: frame_vm_group_bin_4158 (RW)
0x1c3: frame_vm_group_bin_20254 (RW)
0x1c4: frame_vm_group_bin_13058 (RW)
0x1c5: frame_vm_group_bin_5925 (RW)
0x1c6: frame_vm_group_bin_22069 (RW)
0x1c7: frame_vm_group_bin_14917 (RW)
0x1c8: frame_vm_group_bin_7702 (RW)
0x1c9: frame_vm_group_bin_0540 (RW)
0x1c: frame_vm_group_bin_22838 (RW)
0x1ca: frame_vm_group_bin_16732 (RW)
0x1cb: frame_vm_group_bin_9523 (RW)
0x1cc: frame_vm_group_bin_2363 (RW)
0x1cd: frame_vm_group_bin_14810 (RW)
0x1ce: frame_vm_group_bin_11376 (RW)
0x1cf: frame_vm_group_bin_4191 (RW)
0x1d0: frame_vm_group_bin_20286 (RW)
0x1d1: frame_vm_group_bin_13091 (RW)
0x1d2: frame_vm_group_bin_5947 (RW)
0x1d3: frame_vm_group_bin_22099 (RW)
0x1d4: frame_vm_group_bin_14950 (RW)
0x1d5: frame_vm_group_bin_7734 (RW)
0x1d6: frame_vm_group_bin_0571 (RW)
0x1d7: frame_vm_group_bin_16765 (RW)
0x1d8: frame_vm_group_bin_9556 (RW)
0x1d9: frame_vm_group_bin_2396 (RW)
0x1d: frame_vm_group_bin_15655 (RW)
0x1da: frame_vm_group_bin_18491 (RW)
0x1db: frame_vm_group_bin_17979 (RW)
0x1dc: frame_vm_group_bin_4224 (RW)
0x1dd: frame_vm_group_bin_20322 (RW)
0x1de: frame_vm_group_bin_13125 (RW)
0x1df: frame_vm_group_bin_5972 (RW)
0x1e0: frame_vm_group_bin_22133 (RW)
0x1e1: frame_vm_group_bin_14984 (RW)
0x1e2: frame_vm_group_bin_7768 (RW)
0x1e3: frame_vm_group_bin_0604 (RW)
0x1e4: frame_vm_group_bin_16799 (RW)
0x1e5: frame_vm_group_bin_9590 (RW)
0x1e6: frame_vm_group_bin_2429 (RW)
0x1e7: frame_vm_group_bin_18518 (RW)
0x1e8: frame_vm_group_bin_11441 (RW)
0x1e9: frame_vm_group_bin_4257 (RW)
0x1e: frame_vm_group_bin_8465 (RW)
0x1ea: frame_vm_group_bin_20355 (RW)
0x1eb: frame_vm_group_bin_13158 (RW)
0x1ec: frame_vm_group_bin_6003 (RW)
0x1ed: frame_vm_group_bin_22166 (RW)
0x1ee: frame_vm_group_bin_15017 (RW)
0x1ef: frame_vm_group_bin_7801 (RW)
0x1f0: frame_vm_group_bin_0635 (RW)
0x1f1: frame_vm_group_bin_16832 (RW)
0x1f2: frame_vm_group_bin_9623 (RW)
0x1f3: frame_vm_group_bin_2462 (RW)
0x1f4: frame_vm_group_bin_18542 (RW)
0x1f5: frame_vm_group_bin_11474 (RW)
0x1f6: frame_vm_group_bin_4290 (RW)
0x1f7: frame_vm_group_bin_20388 (RW)
0x1f8: frame_vm_group_bin_13191 (RW)
0x1f9: frame_vm_group_bin_6034 (RW)
0x1f: frame_vm_group_bin_1273 (RW)
0x1fa: frame_vm_group_bin_22200 (RW)
0x1fb: frame_vm_group_bin_15046 (RW)
0x1fc: frame_vm_group_bin_7834 (RW)
0x1fd: frame_vm_group_bin_0670 (RW)
0x1fe: frame_vm_group_bin_16865 (RW)
0x1ff: frame_vm_group_bin_9657 (RW)
0x20: frame_vm_group_bin_17469 (RW)
0x21: frame_vm_group_bin_10298 (RW)
0x22: frame_vm_group_bin_3138 (RW)
0x23: frame_vm_group_bin_19207 (RW)
0x24: frame_vm_group_bin_12040 (RW)
0x25: frame_vm_group_bin_4937 (RW)
0x26: frame_vm_group_bin_21032 (RW)
0x27: frame_vm_group_bin_13858 (RW)
0x28: frame_vm_group_bin_6675 (RW)
0x29: frame_vm_group_bin_22871 (RW)
0x2: frame_vm_group_bin_22771 (RW)
0x2a: frame_vm_group_bin_15688 (RW)
0x2b: frame_vm_group_bin_8498 (RW)
0x2c: frame_vm_group_bin_1306 (RW)
0x2d: frame_vm_group_bin_17491 (RW)
0x2e: frame_vm_group_bin_10331 (RW)
0x2f: frame_vm_group_bin_3171 (RW)
0x30: frame_vm_group_bin_19240 (RW)
0x31: frame_vm_group_bin_12067 (RW)
0x32: frame_vm_group_bin_4968 (RW)
0x33: frame_vm_group_bin_21066 (RW)
0x34: frame_vm_group_bin_13888 (RW)
0x35: frame_vm_group_bin_6708 (RW)
0x36: frame_vm_group_bin_22904 (RW)
0x37: frame_vm_group_bin_15721 (RW)
0x38: frame_vm_group_bin_8530 (RW)
0x39: frame_vm_group_bin_1338 (RW)
0x3: frame_vm_group_bin_15588 (RW)
0x3a: frame_vm_group_bin_17517 (RW)
0x3b: frame_vm_group_bin_10365 (RW)
0x3c: frame_vm_group_bin_3205 (RW)
0x3d: frame_vm_group_bin_19274 (RW)
0x3e: frame_vm_group_bin_12101 (RW)
0x3f: frame_vm_group_bin_5002 (RW)
0x40: frame_vm_group_bin_21100 (RW)
0x41: frame_vm_group_bin_13922 (RW)
0x42: frame_vm_group_bin_6741 (RW)
0x43: frame_vm_group_bin_22938 (RW)
0x44: frame_vm_group_bin_15755 (RW)
0x45: frame_vm_group_bin_8562 (RW)
0x46: frame_vm_group_bin_1373 (RW)
0x47: frame_vm_group_bin_17543 (RW)
0x48: frame_vm_group_bin_13193 (RW)
0x49: frame_vm_group_bin_3237 (RW)
0x4: frame_vm_group_bin_8398 (RW)
0x4a: frame_vm_group_bin_19307 (RW)
0x4b: frame_vm_group_bin_12133 (RW)
0x4c: frame_vm_group_bin_5035 (RW)
0x4d: frame_vm_group_bin_21133 (RW)
0x4e: frame_vm_group_bin_13955 (RW)
0x4f: frame_vm_group_bin_6773 (RW)
0x50: frame_vm_group_bin_22970 (RW)
0x51: frame_vm_group_bin_15788 (RW)
0x52: frame_vm_group_bin_8595 (RW)
0x53: frame_vm_group_bin_1406 (RW)
0x54: frame_vm_group_bin_17564 (RW)
0x55: frame_vm_group_bin_10420 (RW)
0x56: frame_vm_group_bin_3270 (RW)
0x57: frame_vm_group_bin_19340 (RW)
0x58: frame_vm_group_bin_12164 (RW)
0x59: frame_vm_group_bin_5069 (RW)
0x5: frame_vm_group_bin_1209 (RW)
0x5a: frame_vm_group_bin_21166 (RW)
0x5b: frame_vm_group_bin_13989 (RW)
0x5c: frame_vm_group_bin_6807 (RW)
0x5d: frame_vm_group_bin_23003 (RW)
0x5e: frame_vm_group_bin_15820 (RW)
0x5f: frame_vm_group_bin_8628 (RW)
0x60: frame_vm_group_bin_1440 (RW)
0x61: frame_vm_group_bin_17589 (RW)
0x62: frame_vm_group_bin_10451 (RW)
0x63: frame_vm_group_bin_3304 (RW)
0x64: frame_vm_group_bin_19374 (RW)
0x65: frame_vm_group_bin_12196 (RW)
0x66: frame_vm_group_bin_5103 (RW)
0x67: frame_vm_group_bin_21199 (RW)
0x68: frame_vm_group_bin_14022 (RW)
0x69: frame_vm_group_bin_12488 (RW)
0x6: frame_vm_group_bin_17423 (RW)
0x6a: frame_vm_group_bin_23036 (RW)
0x6b: frame_vm_group_bin_15853 (RW)
0x6c: frame_vm_group_bin_8661 (RW)
0x6d: frame_vm_group_bin_1473 (RW)
0x6e: frame_vm_group_bin_17613 (RW)
0x6f: frame_vm_group_bin_10484 (RW)
0x70: frame_vm_group_bin_3337 (RW)
0x71: frame_vm_group_bin_19407 (RW)
0x72: frame_vm_group_bin_12226 (RW)
0x73: frame_vm_group_bin_5136 (RW)
0x74: frame_vm_group_bin_21232 (RW)
0x75: frame_vm_group_bin_14055 (RW)
0x76: frame_vm_group_bin_6862 (RW)
0x77: frame_vm_group_bin_23069 (RW)
0x78: frame_vm_group_bin_15886 (RW)
0x79: frame_vm_group_bin_8695 (RW)
0x7: frame_vm_group_bin_10231 (RW)
0x7a: frame_vm_group_bin_1507 (RW)
0x7b: frame_vm_group_bin_17647 (RW)
0x7c: frame_vm_group_bin_10517 (RW)
0x7d: frame_vm_group_bin_3371 (RW)
0x7e: frame_vm_group_bin_19438 (RW)
0x7f: frame_vm_group_bin_12259 (RW)
0x80: frame_vm_group_bin_5170 (RW)
0x81: frame_vm_group_bin_21266 (RW)
0x82: frame_vm_group_bin_14089 (RW)
0x83: frame_vm_group_bin_6888 (RW)
0x84: frame_vm_group_bin_23103 (RW)
0x85: frame_vm_group_bin_15920 (RW)
0x86: frame_vm_group_bin_8729 (RW)
0x87: frame_vm_group_bin_1540 (RW)
0x88: frame_vm_group_bin_17680 (RW)
0x89: frame_vm_group_bin_10550 (RW)
0x8: frame_vm_group_bin_3072 (RW)
0x8a: frame_vm_group_bin_11798 (RW)
0x8b: frame_vm_group_bin_19470 (RW)
0x8c: frame_vm_group_bin_12292 (RW)
0x8d: frame_vm_group_bin_5203 (RW)
0x8e: frame_vm_group_bin_21299 (RW)
0x8f: frame_vm_group_bin_14122 (RW)
0x90: frame_vm_group_bin_6912 (RW)
0x91: frame_vm_group_bin_23136 (RW)
0x92: frame_vm_group_bin_15953 (RW)
0x93: frame_vm_group_bin_8762 (RW)
0x94: frame_vm_group_bin_1573 (RW)
0x95: frame_vm_group_bin_17706 (RW)
0x96: frame_vm_group_bin_10583 (RW)
0x97: frame_vm_group_bin_3423 (RW)
0x98: frame_vm_group_bin_19503 (RW)
0x99: frame_vm_group_bin_12324 (RW)
0x9: frame_vm_group_bin_19140 (RW)
0x9a: frame_vm_group_bin_5237 (RW)
0x9b: frame_vm_group_bin_21331 (RW)
0x9c: frame_vm_group_bin_14156 (RW)
0x9d: frame_vm_group_bin_7855 (RW)
0x9e: frame_vm_group_bin_23169 (RW)
0x9f: frame_vm_group_bin_15989 (RW)
0xa0: frame_vm_group_bin_8796 (RW)
0xa1: frame_vm_group_bin_1607 (RW)
0xa2: frame_vm_group_bin_17734 (RW)
0xa3: frame_vm_group_bin_10617 (RW)
0xa4: frame_vm_group_bin_3446 (RW)
0xa5: frame_vm_group_bin_19537 (RW)
0xa6: frame_vm_group_bin_12358 (RW)
0xa7: frame_vm_group_bin_5270 (RW)
0xa8: frame_vm_group_bin_21364 (RW)
0xa9: frame_vm_group_bin_14188 (RW)
0xa: frame_vm_group_bin_11977 (RW)
0xaa: frame_vm_group_bin_6975 (RW)
0xab: frame_vm_group_bin_11148 (RW)
0xac: frame_vm_group_bin_16022 (RW)
0xad: frame_vm_group_bin_8829 (RW)
0xae: frame_vm_group_bin_1640 (RW)
0xaf: frame_vm_group_bin_17761 (RW)
0xb0: frame_vm_group_bin_10649 (RW)
0xb1: frame_vm_group_bin_3472 (RW)
0xb2: frame_vm_group_bin_19570 (RW)
0xb3: frame_vm_group_bin_12391 (RW)
0xb4: frame_vm_group_bin_5303 (RW)
0xb5: frame_vm_group_bin_21397 (RW)
0xb6: frame_vm_group_bin_14221 (RW)
0xb7: frame_vm_group_bin_7008 (RW)
0xb8: frame_vm_group_bin_23223 (RW)
0xb9: frame_vm_group_bin_16055 (RW)
0xb: frame_vm_group_bin_4872 (RW)
0xba: frame_vm_group_bin_8862 (RW)
0xbb: frame_vm_group_bin_1674 (RW)
0xbc: frame_vm_group_bin_17791 (RW)
0xbd: frame_vm_group_bin_10682 (RW)
0xbe: frame_vm_group_bin_3500 (RW)
0xbf: frame_vm_group_bin_19605 (RW)
0xc0: frame_vm_group_bin_12425 (RW)
0xc1: frame_vm_group_bin_5335 (RW)
0xc2: frame_vm_group_bin_21430 (RW)
0xc3: frame_vm_group_bin_14254 (RW)
0xc4: frame_vm_group_bin_7041 (RW)
0xc5: frame_vm_group_bin_23245 (RW)
0xc6: frame_vm_group_bin_16088 (RW)
0xc7: frame_vm_group_bin_8894 (RW)
0xc8: frame_vm_group_bin_1706 (RW)
0xc9: frame_vm_group_bin_17821 (RW)
0xc: frame_vm_group_bin_20965 (RW)
0xca: frame_vm_group_bin_10714 (RW)
0xcb: frame_vm_group_bin_3528 (RW)
0xcc: frame_vm_group_bin_8671 (RW)
0xcd: frame_vm_group_bin_12456 (RW)
0xce: frame_vm_group_bin_5366 (RW)
0xcf: frame_vm_group_bin_21462 (RW)
0xd0: frame_vm_group_bin_14286 (RW)
0xd1: frame_vm_group_bin_7072 (RW)
0xd2: frame_vm_group_bin_0012 (RW)
0xd3: frame_vm_group_bin_16120 (RW)
0xd4: frame_vm_group_bin_8926 (RW)
0xd5: frame_vm_group_bin_1738 (RW)
0xd6: frame_vm_group_bin_17849 (RW)
0xd7: frame_vm_group_bin_10746 (RW)
0xd8: frame_vm_group_bin_16531 (RW)
0xd9: frame_vm_group_bin_19663 (RW)
0xd: frame_vm_group_bin_13797 (RW)
0xda: frame_vm_group_bin_12489 (RW)
0xdb: frame_vm_group_bin_5399 (RW)
0xdc: frame_vm_group_bin_21494 (RW)
0xdd: frame_vm_group_bin_14318 (RW)
0xde: frame_vm_group_bin_7878 (RW)
0xdf: frame_vm_group_bin_0033 (RW)
0xe0: frame_vm_group_bin_16152 (RW)
0xe1: frame_vm_group_bin_8959 (RW)
0xe2: frame_vm_group_bin_1771 (RW)
0xe3: frame_vm_group_bin_17876 (RW)
0xe4: frame_vm_group_bin_10779 (RW)
0xe5: frame_vm_group_bin_3594 (RW)
0xe6: frame_vm_group_bin_19694 (RW)
0xe7: frame_vm_group_bin_12522 (RW)
0xe8: frame_vm_group_bin_5432 (RW)
0xe9: frame_vm_group_bin_21527 (RW)
0xe: frame_vm_group_bin_6608 (RW)
0xea: frame_vm_group_bin_14351 (RW)
0xeb: frame_vm_group_bin_7136 (RW)
0xec: frame_vm_group_bin_0056 (RW)
0xed: frame_vm_group_bin_16185 (RW)
0xee: frame_vm_group_bin_8992 (RW)
0xef: frame_vm_group_bin_1804 (RW)
0xf0: frame_vm_group_bin_17907 (RW)
0xf1: frame_vm_group_bin_10812 (RW)
0xf2: frame_vm_group_bin_3627 (RW)
0xf3: frame_vm_group_bin_19727 (RW)
0xf4: frame_vm_group_bin_12555 (RW)
0xf5: frame_vm_group_bin_5464 (RW)
0xf6: frame_vm_group_bin_21560 (RW)
0xf7: frame_vm_group_bin_14384 (RW)
0xf8: frame_vm_group_bin_7169 (RW)
0xf9: frame_vm_group_bin_0082 (RW)
0xf: frame_vm_group_bin_22804 (RW)
0xfa: frame_vm_group_bin_16216 (RW)
0xfb: frame_vm_group_bin_9026 (RW)
0xfc: frame_vm_group_bin_1838 (RW)
0xfd: frame_vm_group_bin_17939 (RW)
0xfe: frame_vm_group_bin_10846 (RW)
0xff: frame_vm_group_bin_3661 (RW)
}
pt_vm_group_bin_0026 {
0x0: frame_vm_group_bin_15990 (RW)
0x100: frame_vm_group_bin_21994 (RW)
0x101: frame_vm_group_bin_14818 (RW)
0x102: frame_vm_group_bin_7603 (RW)
0x103: frame_vm_group_bin_0443 (RW)
0x104: frame_vm_group_bin_16633 (RW)
0x105: frame_vm_group_bin_9424 (RW)
0x106: frame_vm_group_bin_2264 (RW)
0x107: frame_vm_group_bin_18367 (RW)
0x108: frame_vm_group_bin_11279 (RW)
0x109: frame_vm_group_bin_4094 (RW)
0x10: frame_vm_group_bin_17762 (RW)
0x10a: frame_vm_group_bin_20188 (RW)
0x10b: frame_vm_group_bin_12990 (RW)
0x10c: frame_vm_group_bin_5873 (RW)
0x10d: frame_vm_group_bin_22023 (RW)
0x10e: frame_vm_group_bin_14851 (RW)
0x10f: frame_vm_group_bin_7636 (RW)
0x110: frame_vm_group_bin_0476 (RW)
0x111: frame_vm_group_bin_16666 (RW)
0x112: frame_vm_group_bin_9457 (RW)
0x113: frame_vm_group_bin_2297 (RW)
0x114: frame_vm_group_bin_18399 (RW)
0x115: frame_vm_group_bin_11312 (RW)
0x116: frame_vm_group_bin_4126 (RW)
0x117: frame_vm_group_bin_20221 (RW)
0x118: frame_vm_group_bin_13025 (RW)
0x119: frame_vm_group_bin_5898 (RW)
0x11: frame_vm_group_bin_10650 (RW)
0x11a: frame_vm_group_bin_22046 (RW)
0x11b: frame_vm_group_bin_14885 (RW)
0x11c: frame_vm_group_bin_7670 (RW)
0x11d: frame_vm_group_bin_0509 (RW)
0x11e: frame_vm_group_bin_16699 (RW)
0x11f: frame_vm_group_bin_9491 (RW)
0x120: frame_vm_group_bin_2331 (RW)
0x121: frame_vm_group_bin_18432 (RW)
0x122: frame_vm_group_bin_11344 (RW)
0x123: frame_vm_group_bin_4159 (RW)
0x124: frame_vm_group_bin_20255 (RW)
0x125: frame_vm_group_bin_13059 (RW)
0x126: frame_vm_group_bin_5926 (RW)
0x127: frame_vm_group_bin_22070 (RW)
0x128: frame_vm_group_bin_14918 (RW)
0x129: frame_vm_group_bin_7703 (RW)
0x12: frame_vm_group_bin_3473 (RW)
0x12a: frame_vm_group_bin_0541 (RW)
0x12b: frame_vm_group_bin_16733 (RW)
0x12c: frame_vm_group_bin_9524 (RW)
0x12d: frame_vm_group_bin_2364 (RW)
0x12e: frame_vm_group_bin_18463 (RW)
0x12f: frame_vm_group_bin_11377 (RW)
0x130: frame_vm_group_bin_4192 (RW)
0x131: frame_vm_group_bin_20287 (RW)
0x132: frame_vm_group_bin_13092 (RW)
0x133: frame_vm_group_bin_5948 (RW)
0x134: frame_vm_group_bin_22100 (RW)
0x135: frame_vm_group_bin_14951 (RW)
0x136: frame_vm_group_bin_7735 (RW)
0x137: frame_vm_group_bin_0572 (RW)
0x138: frame_vm_group_bin_16766 (RW)
0x139: frame_vm_group_bin_9557 (RW)
0x13: frame_vm_group_bin_19571 (RW)
0x13a: frame_vm_group_bin_2398 (RW)
0x13b: frame_vm_group_bin_18492 (RW)
0x13c: frame_vm_group_bin_11409 (RW)
0x13d: frame_vm_group_bin_4225 (RW)
0x13e: frame_vm_group_bin_20323 (RW)
0x13f: frame_vm_group_bin_13126 (RW)
0x140: frame_vm_group_bin_5973 (RW)
0x141: frame_vm_group_bin_22134 (RW)
0x142: frame_vm_group_bin_14985 (RW)
0x143: frame_vm_group_bin_7769 (RW)
0x144: frame_vm_group_bin_0605 (RW)
0x145: frame_vm_group_bin_16800 (RW)
0x146: frame_vm_group_bin_9591 (RW)
0x147: frame_vm_group_bin_2430 (RW)
0x148: frame_vm_group_bin_18519 (RW)
0x149: frame_vm_group_bin_11442 (RW)
0x14: frame_vm_group_bin_12392 (RW)
0x14a: frame_vm_group_bin_4258 (RW)
0x14b: frame_vm_group_bin_20356 (RW)
0x14c: frame_vm_group_bin_13159 (RW)
0x14d: frame_vm_group_bin_6004 (RW)
0x14e: frame_vm_group_bin_22167 (RW)
0x14f: frame_vm_group_bin_15018 (RW)
0x150: frame_vm_group_bin_7802 (RW)
0x151: frame_vm_group_bin_0636 (RW)
0x152: frame_vm_group_bin_16833 (RW)
0x153: frame_vm_group_bin_9624 (RW)
0x154: frame_vm_group_bin_2463 (RW)
0x155: frame_vm_group_bin_18543 (RW)
0x156: frame_vm_group_bin_11475 (RW)
0x157: frame_vm_group_bin_4291 (RW)
0x158: frame_vm_group_bin_20389 (RW)
0x159: frame_vm_group_bin_13192 (RW)
0x15: frame_vm_group_bin_5304 (RW)
0x15a: frame_vm_group_bin_6036 (RW)
0x15b: frame_vm_group_bin_22201 (RW)
0x15c: frame_vm_group_bin_15047 (RW)
0x15d: frame_vm_group_bin_7835 (RW)
0x15e: frame_vm_group_bin_0671 (RW)
0x15f: frame_vm_group_bin_16866 (RW)
0x160: frame_vm_group_bin_9658 (RW)
0x161: frame_vm_group_bin_2496 (RW)
0x162: frame_vm_group_bin_18573 (RW)
0x163: frame_vm_group_bin_11509 (RW)
0x164: frame_vm_group_bin_4325 (RW)
0x165: frame_vm_group_bin_20423 (RW)
0x166: frame_vm_group_bin_13226 (RW)
0x167: frame_vm_group_bin_6061 (RW)
0x168: frame_vm_group_bin_22234 (RW)
0x169: frame_vm_group_bin_15071 (RW)
0x16: frame_vm_group_bin_21398 (RW)
0x16a: frame_vm_group_bin_7868 (RW)
0x16b: frame_vm_group_bin_0704 (RW)
0x16c: frame_vm_group_bin_16898 (RW)
0x16d: frame_vm_group_bin_9690 (RW)
0x16e: frame_vm_group_bin_2529 (RW)
0x16f: frame_vm_group_bin_18606 (RW)
0x170: frame_vm_group_bin_11542 (RW)
0x171: frame_vm_group_bin_4360 (RW)
0x172: frame_vm_group_bin_20456 (RW)
0x173: frame_vm_group_bin_13259 (RW)
0x174: frame_vm_group_bin_6087 (RW)
0x175: frame_vm_group_bin_22267 (RW)
0x176: frame_vm_group_bin_15095 (RW)
0x177: frame_vm_group_bin_7901 (RW)
0x178: frame_vm_group_bin_0737 (RW)
0x179: frame_vm_group_bin_16931 (RW)
0x17: frame_vm_group_bin_14222 (RW)
0x17a: frame_vm_group_bin_9724 (RW)
0x17b: frame_vm_group_bin_2563 (RW)
0x17c: frame_vm_group_bin_18639 (RW)
0x17d: frame_vm_group_bin_11573 (RW)
0x17e: frame_vm_group_bin_4394 (RW)
0x17f: frame_vm_group_bin_20490 (RW)
0x180: frame_vm_group_bin_13293 (RW)
0x181: frame_vm_group_bin_6118 (RW)
0x182: frame_vm_group_bin_22300 (RW)
0x183: frame_vm_group_bin_15125 (RW)
0x184: frame_vm_group_bin_7936 (RW)
0x185: frame_vm_group_bin_0771 (RW)
0x186: frame_vm_group_bin_16965 (RW)
0x187: frame_vm_group_bin_9757 (RW)
0x188: frame_vm_group_bin_2596 (RW)
0x189: frame_vm_group_bin_18672 (RW)
0x18: frame_vm_group_bin_7009 (RW)
0x18a: frame_vm_group_bin_11598 (RW)
0x18b: frame_vm_group_bin_4427 (RW)
0x18c: frame_vm_group_bin_20523 (RW)
0x18d: frame_vm_group_bin_13325 (RW)
0x18e: frame_vm_group_bin_6150 (RW)
0x18f: frame_vm_group_bin_22333 (RW)
0x190: frame_vm_group_bin_15148 (RW)
0x191: frame_vm_group_bin_7969 (RW)
0x192: frame_vm_group_bin_0804 (RW)
0x193: frame_vm_group_bin_16998 (RW)
0x194: frame_vm_group_bin_9790 (RW)
0x195: frame_vm_group_bin_2629 (RW)
0x196: frame_vm_group_bin_18704 (RW)
0x197: frame_vm_group_bin_11623 (RW)
0x198: frame_vm_group_bin_4460 (RW)
0x199: frame_vm_group_bin_20556 (RW)
0x19: frame_vm_group_bin_23224 (RW)
0x19a: frame_vm_group_bin_13359 (RW)
0x19b: frame_vm_group_bin_6184 (RW)
0x19c: frame_vm_group_bin_22366 (RW)
0x19d: frame_vm_group_bin_15182 (RW)
0x19e: frame_vm_group_bin_8001 (RW)
0x19f: frame_vm_group_bin_0837 (RW)
0x1: frame_vm_group_bin_8797 (RW)
0x1a0: frame_vm_group_bin_17032 (RW)
0x1a1: frame_vm_group_bin_9824 (RW)
0x1a2: frame_vm_group_bin_2663 (RW)
0x1a3: frame_vm_group_bin_18736 (RW)
0x1a4: frame_vm_group_bin_11647 (RW)
0x1a5: frame_vm_group_bin_4494 (RW)
0x1a6: frame_vm_group_bin_20590 (RW)
0x1a7: frame_vm_group_bin_13390 (RW)
0x1a8: frame_vm_group_bin_6212 (RW)
0x1a9: frame_vm_group_bin_22399 (RW)
0x1a: frame_vm_group_bin_16057 (RW)
0x1aa: frame_vm_group_bin_15215 (RW)
0x1ab: frame_vm_group_bin_8029 (RW)
0x1ac: frame_vm_group_bin_0870 (RW)
0x1ad: frame_vm_group_bin_17065 (RW)
0x1ae: frame_vm_group_bin_9857 (RW)
0x1af: frame_vm_group_bin_2696 (RW)
0x1b0: frame_vm_group_bin_18769 (RW)
0x1b1: frame_vm_group_bin_11668 (RW)
0x1b2: frame_vm_group_bin_4527 (RW)
0x1b3: frame_vm_group_bin_20623 (RW)
0x1b4: frame_vm_group_bin_13423 (RW)
0x1b5: frame_vm_group_bin_6240 (RW)
0x1b6: frame_vm_group_bin_22431 (RW)
0x1b7: frame_vm_group_bin_15249 (RW)
0x1b8: frame_vm_group_bin_8059 (RW)
0x1b9: frame_vm_group_bin_0903 (RW)
0x1b: frame_vm_group_bin_8863 (RW)
0x1ba: frame_vm_group_bin_17099 (RW)
0x1bb: frame_vm_group_bin_9890 (RW)
0x1bc: frame_vm_group_bin_2730 (RW)
0x1bd: frame_vm_group_bin_18803 (RW)
0x1be: frame_vm_group_bin_11695 (RW)
0x1bf: frame_vm_group_bin_4560 (RW)
0x1c0: frame_vm_group_bin_20656 (RW)
0x1c1: frame_vm_group_bin_13457 (RW)
0x1c2: frame_vm_group_bin_6272 (RW)
0x1c3: frame_vm_group_bin_22465 (RW)
0x1c4: frame_vm_group_bin_15282 (RW)
0x1c5: frame_vm_group_bin_8092 (RW)
0x1c6: frame_vm_group_bin_0937 (RW)
0x1c7: frame_vm_group_bin_17132 (RW)
0x1c8: frame_vm_group_bin_9923 (RW)
0x1c9: frame_vm_group_bin_2763 (RW)
0x1c: frame_vm_group_bin_1675 (RW)
0x1ca: frame_vm_group_bin_18837 (RW)
0x1cb: frame_vm_group_bin_11723 (RW)
0x1cc: frame_vm_group_bin_4585 (RW)
0x1cd: frame_vm_group_bin_20689 (RW)
0x1ce: frame_vm_group_bin_13490 (RW)
0x1cf: frame_vm_group_bin_6305 (RW)
0x1d0: frame_vm_group_bin_22498 (RW)
0x1d1: frame_vm_group_bin_15315 (RW)
0x1d2: frame_vm_group_bin_8124 (RW)
0x1d3: frame_vm_group_bin_0970 (RW)
0x1d4: frame_vm_group_bin_17164 (RW)
0x1d5: frame_vm_group_bin_9954 (RW)
0x1d6: frame_vm_group_bin_2796 (RW)
0x1d7: frame_vm_group_bin_18870 (RW)
0x1d8: frame_vm_group_bin_11745 (RW)
0x1d9: frame_vm_group_bin_4608 (RW)
0x1d: frame_vm_group_bin_17792 (RW)
0x1da: frame_vm_group_bin_20723 (RW)
0x1db: frame_vm_group_bin_13524 (RW)
0x1dc: frame_vm_group_bin_6338 (RW)
0x1dd: frame_vm_group_bin_22531 (RW)
0x1de: frame_vm_group_bin_15349 (RW)
0x1df: frame_vm_group_bin_8158 (RW)
0x1e0: frame_vm_group_bin_1004 (RW)
0x1e1: frame_vm_group_bin_17195 (RW)
0x1e2: frame_vm_group_bin_9988 (RW)
0x1e3: frame_vm_group_bin_2830 (RW)
0x1e4: frame_vm_group_bin_18904 (RW)
0x1e5: frame_vm_group_bin_11769 (RW)
0x1e6: frame_vm_group_bin_4635 (RW)
0x1e7: frame_vm_group_bin_20756 (RW)
0x1e8: frame_vm_group_bin_13557 (RW)
0x1e9: frame_vm_group_bin_6371 (RW)
0x1e: frame_vm_group_bin_10683 (RW)
0x1ea: frame_vm_group_bin_22564 (RW)
0x1eb: frame_vm_group_bin_15382 (RW)
0x1ec: frame_vm_group_bin_8191 (RW)
0x1ed: frame_vm_group_bin_1029 (RW)
0x1ee: frame_vm_group_bin_17228 (RW)
0x1ef: frame_vm_group_bin_10021 (RW)
0x1f0: frame_vm_group_bin_2862 (RW)
0x1f1: frame_vm_group_bin_18937 (RW)
0x1f2: frame_vm_group_bin_11794 (RW)
0x1f3: frame_vm_group_bin_4668 (RW)
0x1f4: frame_vm_group_bin_20789 (RW)
0x1f5: frame_vm_group_bin_13590 (RW)
0x1f6: frame_vm_group_bin_6401 (RW)
0x1f7: frame_vm_group_bin_22597 (RW)
0x1f8: frame_vm_group_bin_15415 (RW)
0x1f9: frame_vm_group_bin_8224 (RW)
0x1f: frame_vm_group_bin_3501 (RW)
0x1fa: frame_vm_group_bin_1052 (RW)
0x1fb: frame_vm_group_bin_17261 (RW)
0x1fc: frame_vm_group_bin_10055 (RW)
0x1fd: frame_vm_group_bin_2898 (RW)
0x1fe: frame_vm_group_bin_18969 (RW)
0x1ff: frame_vm_group_bin_11827 (RW)
0x20: frame_vm_group_bin_19606 (RW)
0x21: frame_vm_group_bin_12426 (RW)
0x22: frame_vm_group_bin_5336 (RW)
0x23: frame_vm_group_bin_21431 (RW)
0x24: frame_vm_group_bin_14255 (RW)
0x25: frame_vm_group_bin_7042 (RW)
0x26: frame_vm_group_bin_23246 (RW)
0x27: frame_vm_group_bin_16089 (RW)
0x28: frame_vm_group_bin_8895 (RW)
0x29: frame_vm_group_bin_1707 (RW)
0x2: frame_vm_group_bin_1608 (RW)
0x2a: frame_vm_group_bin_17822 (RW)
0x2b: frame_vm_group_bin_10715 (RW)
0x2c: frame_vm_group_bin_3529 (RW)
0x2d: frame_vm_group_bin_19637 (RW)
0x2e: frame_vm_group_bin_12457 (RW)
0x2f: frame_vm_group_bin_5367 (RW)
0x30: frame_vm_group_bin_21463 (RW)
0x31: frame_vm_group_bin_14287 (RW)
0x32: frame_vm_group_bin_7073 (RW)
0x33: frame_vm_group_bin_0013 (RW)
0x34: frame_vm_group_bin_16121 (RW)
0x35: frame_vm_group_bin_8927 (RW)
0x36: frame_vm_group_bin_1739 (RW)
0x37: frame_vm_group_bin_17850 (RW)
0x38: frame_vm_group_bin_10747 (RW)
0x39: frame_vm_group_bin_3560 (RW)
0x3: frame_vm_group_bin_17735 (RW)
0x3a: frame_vm_group_bin_19665 (RW)
0x3b: frame_vm_group_bin_12490 (RW)
0x3c: frame_vm_group_bin_5400 (RW)
0x3d: frame_vm_group_bin_21495 (RW)
0x3e: frame_vm_group_bin_14319 (RW)
0x3f: frame_vm_group_bin_7105 (RW)
0x40: frame_vm_group_bin_0034 (RW)
0x41: frame_vm_group_bin_16153 (RW)
0x42: frame_vm_group_bin_8960 (RW)
0x43: frame_vm_group_bin_1772 (RW)
0x44: frame_vm_group_bin_17877 (RW)
0x45: frame_vm_group_bin_10780 (RW)
0x46: frame_vm_group_bin_3595 (RW)
0x47: frame_vm_group_bin_19695 (RW)
0x48: frame_vm_group_bin_12523 (RW)
0x49: frame_vm_group_bin_5433 (RW)
0x4: frame_vm_group_bin_10618 (RW)
0x4a: frame_vm_group_bin_21528 (RW)
0x4b: frame_vm_group_bin_14352 (RW)
0x4c: frame_vm_group_bin_7137 (RW)
0x4d: frame_vm_group_bin_0057 (RW)
0x4e: frame_vm_group_bin_16186 (RW)
0x4f: frame_vm_group_bin_8993 (RW)
0x50: frame_vm_group_bin_1805 (RW)
0x51: frame_vm_group_bin_17908 (RW)
0x52: frame_vm_group_bin_10813 (RW)
0x53: frame_vm_group_bin_3628 (RW)
0x54: frame_vm_group_bin_19728 (RW)
0x55: frame_vm_group_bin_12556 (RW)
0x56: frame_vm_group_bin_5465 (RW)
0x57: frame_vm_group_bin_21561 (RW)
0x58: frame_vm_group_bin_14385 (RW)
0x59: frame_vm_group_bin_7172 (RW)
0x5: frame_vm_group_bin_3447 (RW)
0x5a: frame_vm_group_bin_0084 (RW)
0x5b: frame_vm_group_bin_16217 (RW)
0x5c: frame_vm_group_bin_9027 (RW)
0x5d: frame_vm_group_bin_1839 (RW)
0x5e: frame_vm_group_bin_17940 (RW)
0x5f: frame_vm_group_bin_10847 (RW)
0x60: frame_vm_group_bin_3662 (RW)
0x61: frame_vm_group_bin_19762 (RW)
0x62: frame_vm_group_bin_12590 (RW)
0x63: frame_vm_group_bin_5498 (RW)
0x64: frame_vm_group_bin_21595 (RW)
0x65: frame_vm_group_bin_14419 (RW)
0x66: frame_vm_group_bin_7206 (RW)
0x67: frame_vm_group_bin_0109 (RW)
0x68: frame_vm_group_bin_16243 (RW)
0x69: frame_vm_group_bin_9060 (RW)
0x6: frame_vm_group_bin_19538 (RW)
0x6a: frame_vm_group_bin_1872 (RW)
0x6b: frame_vm_group_bin_17972 (RW)
0x6c: frame_vm_group_bin_10879 (RW)
0x6d: frame_vm_group_bin_3695 (RW)
0x6e: frame_vm_group_bin_19795 (RW)
0x6f: frame_vm_group_bin_12623 (RW)
0x70: frame_vm_group_bin_5530 (RW)
0x71: frame_vm_group_bin_21628 (RW)
0x72: frame_vm_group_bin_14452 (RW)
0x73: frame_vm_group_bin_7239 (RW)
0x74: frame_vm_group_bin_0131 (RW)
0x75: frame_vm_group_bin_16270 (RW)
0x76: frame_vm_group_bin_9093 (RW)
0x77: frame_vm_group_bin_1905 (RW)
0x78: frame_vm_group_bin_18003 (RW)
0x79: frame_vm_group_bin_10913 (RW)
0x7: frame_vm_group_bin_12359 (RW)
0x7a: frame_vm_group_bin_3729 (RW)
0x7b: frame_vm_group_bin_19829 (RW)
0x7c: frame_vm_group_bin_12655 (RW)
0x7d: frame_vm_group_bin_5564 (RW)
0x7e: frame_vm_group_bin_21662 (RW)
0x7f: frame_vm_group_bin_14486 (RW)
0x80: frame_vm_group_bin_7273 (RW)
0x81: frame_vm_group_bin_0154 (RW)
0x82: frame_vm_group_bin_16302 (RW)
0x83: frame_vm_group_bin_9127 (RW)
0x84: frame_vm_group_bin_1939 (RW)
0x85: frame_vm_group_bin_18037 (RW)
0x86: frame_vm_group_bin_10947 (RW)
0x87: frame_vm_group_bin_3762 (RW)
0x88: frame_vm_group_bin_19862 (RW)
0x89: frame_vm_group_bin_12679 (RW)
0x8: frame_vm_group_bin_5271 (RW)
0x8a: frame_vm_group_bin_5596 (RW)
0x8b: frame_vm_group_bin_21694 (RW)
0x8c: frame_vm_group_bin_14520 (RW)
0x8d: frame_vm_group_bin_7305 (RW)
0x8e: frame_vm_group_bin_0180 (RW)
0x8f: frame_vm_group_bin_16334 (RW)
0x90: frame_vm_group_bin_9159 (RW)
0x91: frame_vm_group_bin_1971 (RW)
0x92: frame_vm_group_bin_18069 (RW)
0x93: frame_vm_group_bin_10979 (RW)
0x94: frame_vm_group_bin_3794 (RW)
0x95: frame_vm_group_bin_19894 (RW)
0x96: frame_vm_group_bin_12703 (RW)
0x97: frame_vm_group_bin_5627 (RW)
0x98: frame_vm_group_bin_21727 (RW)
0x99: frame_vm_group_bin_14553 (RW)
0x9: frame_vm_group_bin_21365 (RW)
0x9a: frame_vm_group_bin_7339 (RW)
0x9b: frame_vm_group_bin_0213 (RW)
0x9c: frame_vm_group_bin_16368 (RW)
0x9d: frame_vm_group_bin_9191 (RW)
0x9e: frame_vm_group_bin_2005 (RW)
0x9f: frame_vm_group_bin_18101 (RW)
0xa0: frame_vm_group_bin_11013 (RW)
0xa1: frame_vm_group_bin_3828 (RW)
0xa2: frame_vm_group_bin_19926 (RW)
0xa3: frame_vm_group_bin_12730 (RW)
0xa4: frame_vm_group_bin_5661 (RW)
0xa5: frame_vm_group_bin_21761 (RW)
0xa6: frame_vm_group_bin_14587 (RW)
0xa7: frame_vm_group_bin_7372 (RW)
0xa8: frame_vm_group_bin_0240 (RW)
0xa9: frame_vm_group_bin_16401 (RW)
0xa: frame_vm_group_bin_14189 (RW)
0xaa: frame_vm_group_bin_9218 (RW)
0xab: frame_vm_group_bin_2038 (RW)
0xac: frame_vm_group_bin_18134 (RW)
0xad: frame_vm_group_bin_11046 (RW)
0xae: frame_vm_group_bin_3861 (RW)
0xaf: frame_vm_group_bin_19959 (RW)
0xb0: frame_vm_group_bin_12758 (RW)
0xb1: frame_vm_group_bin_5694 (RW)
0xb2: frame_vm_group_bin_21793 (RW)
0xb3: frame_vm_group_bin_14619 (RW)
0xb4: frame_vm_group_bin_7405 (RW)
0xb5: frame_vm_group_bin_0261 (RW)
0xb6: frame_vm_group_bin_16434 (RW)
0xb7: frame_vm_group_bin_9242 (RW)
0xb8: frame_vm_group_bin_2071 (RW)
0xb9: frame_vm_group_bin_18167 (RW)
0xb: frame_vm_group_bin_6976 (RW)
0xba: frame_vm_group_bin_11080 (RW)
0xbb: frame_vm_group_bin_3895 (RW)
0xbc: frame_vm_group_bin_19991 (RW)
0xbd: frame_vm_group_bin_12792 (RW)
0xbe: frame_vm_group_bin_5728 (RW)
0xbf: frame_vm_group_bin_21828 (RW)
0xc0: frame_vm_group_bin_14653 (RW)
0xc1: frame_vm_group_bin_7439 (RW)
0xc2: frame_vm_group_bin_0288 (RW)
0xc3: frame_vm_group_bin_16468 (RW)
0xc4: frame_vm_group_bin_9266 (RW)
0xc5: frame_vm_group_bin_2105 (RW)
0xc6: frame_vm_group_bin_18200 (RW)
0xc7: frame_vm_group_bin_11113 (RW)
0xc8: frame_vm_group_bin_3928 (RW)
0xc9: frame_vm_group_bin_20024 (RW)
0xc: frame_vm_group_bin_23201 (RW)
0xca: frame_vm_group_bin_12824 (RW)
0xcb: frame_vm_group_bin_5754 (RW)
0xcc: frame_vm_group_bin_21861 (RW)
0xcd: frame_vm_group_bin_14686 (RW)
0xce: frame_vm_group_bin_7472 (RW)
0xcf: frame_vm_group_bin_0319 (RW)
0xd0: frame_vm_group_bin_16501 (RW)
0xd1: frame_vm_group_bin_9292 (RW)
0xd2: frame_vm_group_bin_2139 (RW)
0xd3: frame_vm_group_bin_18233 (RW)
0xd4: frame_vm_group_bin_11145 (RW)
0xd5: frame_vm_group_bin_3960 (RW)
0xd6: frame_vm_group_bin_20057 (RW)
0xd7: frame_vm_group_bin_12857 (RW)
0xd8: frame_vm_group_bin_5778 (RW)
0xd9: frame_vm_group_bin_21894 (RW)
0xd: frame_vm_group_bin_16023 (RW)
0xda: frame_vm_group_bin_14720 (RW)
0xdb: frame_vm_group_bin_7505 (RW)
0xdc: frame_vm_group_bin_0351 (RW)
0xdd: frame_vm_group_bin_16535 (RW)
0xde: frame_vm_group_bin_9323 (RW)
0xdf: frame_vm_group_bin_2173 (RW)
0xe0: frame_vm_group_bin_18267 (RW)
0xe1: frame_vm_group_bin_11179 (RW)
0xe2: frame_vm_group_bin_3994 (RW)
0xe3: frame_vm_group_bin_20091 (RW)
0xe4: frame_vm_group_bin_12891 (RW)
0xe5: frame_vm_group_bin_5801 (RW)
0xe6: frame_vm_group_bin_21927 (RW)
0xe7: frame_vm_group_bin_14752 (RW)
0xe8: frame_vm_group_bin_7537 (RW)
0xe9: frame_vm_group_bin_0383 (RW)
0xe: frame_vm_group_bin_8830 (RW)
0xea: frame_vm_group_bin_16567 (RW)
0xeb: frame_vm_group_bin_9356 (RW)
0xec: frame_vm_group_bin_2204 (RW)
0xed: frame_vm_group_bin_18300 (RW)
0xee: frame_vm_group_bin_11212 (RW)
0xef: frame_vm_group_bin_4027 (RW)
0xf0: frame_vm_group_bin_20123 (RW)
0xf1: frame_vm_group_bin_12924 (RW)
0xf2: frame_vm_group_bin_5822 (RW)
0xf3: frame_vm_group_bin_21960 (RW)
0xf4: frame_vm_group_bin_14784 (RW)
0xf5: frame_vm_group_bin_7569 (RW)
0xf6: frame_vm_group_bin_0411 (RW)
0xf7: frame_vm_group_bin_16599 (RW)
0xf8: frame_vm_group_bin_9389 (RW)
0xf9: frame_vm_group_bin_2232 (RW)
0xf: frame_vm_group_bin_1641 (RW)
0xfa: frame_vm_group_bin_18334 (RW)
0xfb: frame_vm_group_bin_11246 (RW)
0xfc: frame_vm_group_bin_4061 (RW)
0xfd: frame_vm_group_bin_20156 (RW)
0xfe: frame_vm_group_bin_12957 (RW)
0xff: frame_vm_group_bin_5848 (RW)
}
pt_vm_group_bin_0028 {
0x0: frame_vm_group_bin_0647 (RW)
0x100: frame_vm_group_bin_6644 (RW)
0x101: frame_vm_group_bin_22840 (RW)
0x102: frame_vm_group_bin_15657 (RW)
0x103: frame_vm_group_bin_8467 (RW)
0x104: frame_vm_group_bin_1275 (RW)
0x105: frame_vm_group_bin_17471 (RW)
0x106: frame_vm_group_bin_10300 (RW)
0x107: frame_vm_group_bin_3140 (RW)
0x108: frame_vm_group_bin_19209 (RW)
0x109: frame_vm_group_bin_12042 (RW)
0x10: frame_vm_group_bin_2505 (RW)
0x10a: frame_vm_group_bin_4939 (RW)
0x10b: frame_vm_group_bin_21034 (RW)
0x10c: frame_vm_group_bin_13860 (RW)
0x10d: frame_vm_group_bin_6677 (RW)
0x10e: frame_vm_group_bin_22873 (RW)
0x10f: frame_vm_group_bin_15690 (RW)
0x110: frame_vm_group_bin_8500 (RW)
0x111: frame_vm_group_bin_1308 (RW)
0x112: frame_vm_group_bin_17493 (RW)
0x113: frame_vm_group_bin_10333 (RW)
0x114: frame_vm_group_bin_3173 (RW)
0x115: frame_vm_group_bin_19242 (RW)
0x116: frame_vm_group_bin_12069 (RW)
0x117: frame_vm_group_bin_4970 (RW)
0x118: frame_vm_group_bin_21068 (RW)
0x119: frame_vm_group_bin_13890 (RW)
0x11: frame_vm_group_bin_18582 (RW)
0x11a: frame_vm_group_bin_6711 (RW)
0x11b: frame_vm_group_bin_22907 (RW)
0x11c: frame_vm_group_bin_15724 (RW)
0x11d: frame_vm_group_bin_8533 (RW)
0x11e: frame_vm_group_bin_1341 (RW)
0x11f: frame_vm_group_bin_17519 (RW)
0x120: frame_vm_group_bin_10367 (RW)
0x121: frame_vm_group_bin_3207 (RW)
0x122: frame_vm_group_bin_19276 (RW)
0x123: frame_vm_group_bin_12103 (RW)
0x124: frame_vm_group_bin_5004 (RW)
0x125: frame_vm_group_bin_21102 (RW)
0x126: frame_vm_group_bin_13924 (RW)
0x127: frame_vm_group_bin_6743 (RW)
0x128: frame_vm_group_bin_22940 (RW)
0x129: frame_vm_group_bin_15757 (RW)
0x12: frame_vm_group_bin_11518 (RW)
0x12a: frame_vm_group_bin_8564 (RW)
0x12b: frame_vm_group_bin_1375 (RW)
0x12c: frame_vm_group_bin_12558 (RW)
0x12d: frame_vm_group_bin_10396 (RW)
0x12e: frame_vm_group_bin_3239 (RW)
0x12f: frame_vm_group_bin_19309 (RW)
0x130: frame_vm_group_bin_12135 (RW)
0x131: frame_vm_group_bin_5037 (RW)
0x132: frame_vm_group_bin_21135 (RW)
0x133: frame_vm_group_bin_13957 (RW)
0x134: frame_vm_group_bin_6775 (RW)
0x135: frame_vm_group_bin_22972 (RW)
0x136: frame_vm_group_bin_15790 (RW)
0x137: frame_vm_group_bin_8597 (RW)
0x138: frame_vm_group_bin_1408 (RW)
0x139: frame_vm_group_bin_17566 (RW)
0x13: frame_vm_group_bin_4334 (RW)
0x13a: frame_vm_group_bin_10423 (RW)
0x13b: frame_vm_group_bin_3273 (RW)
0x13c: frame_vm_group_bin_19343 (RW)
0x13d: frame_vm_group_bin_11569 (RW)
0x13e: frame_vm_group_bin_5072 (RW)
0x13f: frame_vm_group_bin_21168 (RW)
0x140: frame_vm_group_bin_13991 (RW)
0x141: frame_vm_group_bin_5810 (RW)
0x142: frame_vm_group_bin_23005 (RW)
0x143: frame_vm_group_bin_15822 (RW)
0x144: frame_vm_group_bin_8630 (RW)
0x145: frame_vm_group_bin_1442 (RW)
0x146: frame_vm_group_bin_21941 (RW)
0x147: frame_vm_group_bin_10453 (RW)
0x148: frame_vm_group_bin_3306 (RW)
0x149: frame_vm_group_bin_19376 (RW)
0x14: frame_vm_group_bin_20432 (RW)
0x14a: frame_vm_group_bin_12198 (RW)
0x14b: frame_vm_group_bin_5105 (RW)
0x14c: frame_vm_group_bin_21201 (RW)
0x14d: frame_vm_group_bin_14024 (RW)
0x14e: frame_vm_group_bin_6837 (RW)
0x14f: frame_vm_group_bin_23038 (RW)
0x150: frame_vm_group_bin_15855 (RW)
0x151: frame_vm_group_bin_8663 (RW)
0x152: frame_vm_group_bin_1475 (RW)
0x153: frame_vm_group_bin_17615 (RW)
0x154: frame_vm_group_bin_10486 (RW)
0x155: frame_vm_group_bin_3339 (RW)
0x156: frame_vm_group_bin_19409 (RW)
0x157: frame_vm_group_bin_12228 (RW)
0x158: frame_vm_group_bin_5138 (RW)
0x159: frame_vm_group_bin_21234 (RW)
0x15: frame_vm_group_bin_13235 (RW)
0x15a: frame_vm_group_bin_14058 (RW)
0x15b: frame_vm_group_bin_6865 (RW)
0x15c: frame_vm_group_bin_23072 (RW)
0x15d: frame_vm_group_bin_15889 (RW)
0x15e: frame_vm_group_bin_8698 (RW)
0x15f: frame_vm_group_bin_1509 (RW)
0x160: frame_vm_group_bin_17649 (RW)
0x161: frame_vm_group_bin_10519 (RW)
0x162: frame_vm_group_bin_3373 (RW)
0x163: frame_vm_group_bin_19440 (RW)
0x164: frame_vm_group_bin_12261 (RW)
0x165: frame_vm_group_bin_5172 (RW)
0x166: frame_vm_group_bin_21268 (RW)
0x167: frame_vm_group_bin_14091 (RW)
0x168: frame_vm_group_bin_6890 (RW)
0x169: frame_vm_group_bin_23105 (RW)
0x16: frame_vm_group_bin_15026 (RW)
0x16a: frame_vm_group_bin_15922 (RW)
0x16b: frame_vm_group_bin_8731 (RW)
0x16c: frame_vm_group_bin_1542 (RW)
0x16d: frame_vm_group_bin_12582 (RW)
0x16e: frame_vm_group_bin_10552 (RW)
0x16f: frame_vm_group_bin_3401 (RW)
0x170: frame_vm_group_bin_19472 (RW)
0x171: frame_vm_group_bin_12294 (RW)
0x172: frame_vm_group_bin_5205 (RW)
0x173: frame_vm_group_bin_21301 (RW)
0x174: frame_vm_group_bin_14124 (RW)
0x175: frame_vm_group_bin_6914 (RW)
0x176: frame_vm_group_bin_23138 (RW)
0x177: frame_vm_group_bin_15955 (RW)
0x178: frame_vm_group_bin_8764 (RW)
0x179: frame_vm_group_bin_1575 (RW)
0x17: frame_vm_group_bin_22243 (RW)
0x17a: frame_vm_group_bin_17709 (RW)
0x17b: frame_vm_group_bin_10586 (RW)
0x17c: frame_vm_group_bin_3426 (RW)
0x17d: frame_vm_group_bin_19506 (RW)
0x17e: frame_vm_group_bin_12327 (RW)
0x17f: frame_vm_group_bin_5239 (RW)
0x180: frame_vm_group_bin_21333 (RW)
0x181: frame_vm_group_bin_14158 (RW)
0x182: frame_vm_group_bin_6945 (RW)
0x183: frame_vm_group_bin_23171 (RW)
0x184: frame_vm_group_bin_15991 (RW)
0x185: frame_vm_group_bin_8798 (RW)
0x186: frame_vm_group_bin_1609 (RW)
0x187: frame_vm_group_bin_21964 (RW)
0x188: frame_vm_group_bin_10619 (RW)
0x189: frame_vm_group_bin_3448 (RW)
0x18: frame_vm_group_bin_15077 (RW)
0x18a: frame_vm_group_bin_19539 (RW)
0x18b: frame_vm_group_bin_12360 (RW)
0x18c: frame_vm_group_bin_5272 (RW)
0x18d: frame_vm_group_bin_21366 (RW)
0x18e: frame_vm_group_bin_14190 (RW)
0x18f: frame_vm_group_bin_6977 (RW)
0x190: frame_vm_group_bin_23202 (RW)
0x191: frame_vm_group_bin_16024 (RW)
0x192: frame_vm_group_bin_8831 (RW)
0x193: frame_vm_group_bin_1642 (RW)
0x194: frame_vm_group_bin_3344 (RW)
0x195: frame_vm_group_bin_10651 (RW)
0x196: frame_vm_group_bin_3474 (RW)
0x197: frame_vm_group_bin_19572 (RW)
0x198: frame_vm_group_bin_12393 (RW)
0x199: frame_vm_group_bin_5305 (RW)
0x19: frame_vm_group_bin_7877 (RW)
0x19a: frame_vm_group_bin_21400 (RW)
0x19b: frame_vm_group_bin_14224 (RW)
0x19c: frame_vm_group_bin_7011 (RW)
0x19d: frame_vm_group_bin_23226 (RW)
0x19e: frame_vm_group_bin_16058 (RW)
0x19f: frame_vm_group_bin_8864 (RW)
0x1: frame_vm_group_bin_16843 (RW)
0x1a0: frame_vm_group_bin_1676 (RW)
0x1a1: frame_vm_group_bin_17793 (RW)
0x1a2: frame_vm_group_bin_10684 (RW)
0x1a3: frame_vm_group_bin_3502 (RW)
0x1a4: frame_vm_group_bin_19607 (RW)
0x1a5: frame_vm_group_bin_12427 (RW)
0x1a6: frame_vm_group_bin_5337 (RW)
0x1a7: frame_vm_group_bin_21432 (RW)
0x1a8: frame_vm_group_bin_14256 (RW)
0x1a9: frame_vm_group_bin_7043 (RW)
0x1a: frame_vm_group_bin_0714 (RW)
0x1aa: frame_vm_group_bin_23247 (RW)
0x1ab: frame_vm_group_bin_16090 (RW)
0x1ac: frame_vm_group_bin_8896 (RW)
0x1ad: frame_vm_group_bin_1708 (RW)
0x1ae: frame_vm_group_bin_17823 (RW)
0x1af: frame_vm_group_bin_10716 (RW)
0x1b0: frame_vm_group_bin_3530 (RW)
0x1b1: frame_vm_group_bin_19638 (RW)
0x1b2: frame_vm_group_bin_12458 (RW)
0x1b3: frame_vm_group_bin_5368 (RW)
0x1b4: frame_vm_group_bin_21464 (RW)
0x1b5: frame_vm_group_bin_14288 (RW)
0x1b6: frame_vm_group_bin_7074 (RW)
0x1b7: frame_vm_group_bin_0014 (RW)
0x1b8: frame_vm_group_bin_16122 (RW)
0x1b9: frame_vm_group_bin_8928 (RW)
0x1b: frame_vm_group_bin_16908 (RW)
0x1ba: frame_vm_group_bin_1741 (RW)
0x1bb: frame_vm_group_bin_17852 (RW)
0x1bc: frame_vm_group_bin_10749 (RW)
0x1bd: frame_vm_group_bin_3562 (RW)
0x1be: frame_vm_group_bin_19666 (RW)
0x1bf: frame_vm_group_bin_12491 (RW)
0x1c0: frame_vm_group_bin_5401 (RW)
0x1c1: frame_vm_group_bin_21496 (RW)
0x1c2: frame_vm_group_bin_14320 (RW)
0x1c3: frame_vm_group_bin_7106 (RW)
0x1c4: frame_vm_group_bin_4436 (RW)
0x1c5: frame_vm_group_bin_16154 (RW)
0x1c6: frame_vm_group_bin_8961 (RW)
0x1c7: frame_vm_group_bin_1773 (RW)
0x1c8: frame_vm_group_bin_21987 (RW)
0x1c9: frame_vm_group_bin_10781 (RW)
0x1c: frame_vm_group_bin_9700 (RW)
0x1ca: frame_vm_group_bin_3596 (RW)
0x1cb: frame_vm_group_bin_19696 (RW)
0x1cc: frame_vm_group_bin_12524 (RW)
0x1cd: frame_vm_group_bin_5434 (RW)
0x1ce: frame_vm_group_bin_21529 (RW)
0x1cf: frame_vm_group_bin_14353 (RW)
0x1d0: frame_vm_group_bin_7138 (RW)
0x1d1: frame_vm_group_bin_9071 (RW)
0x1d2: frame_vm_group_bin_16187 (RW)
0x1d3: frame_vm_group_bin_8994 (RW)
0x1d4: frame_vm_group_bin_1806 (RW)
0x1d5: frame_vm_group_bin_17909 (RW)
0x1d6: frame_vm_group_bin_10814 (RW)
0x1d7: frame_vm_group_bin_3629 (RW)
0x1d8: frame_vm_group_bin_19729 (RW)
0x1d9: frame_vm_group_bin_12557 (RW)
0x1d: frame_vm_group_bin_2539 (RW)
0x1da: frame_vm_group_bin_5467 (RW)
0x1db: frame_vm_group_bin_21563 (RW)
0x1dc: frame_vm_group_bin_14387 (RW)
0x1dd: frame_vm_group_bin_7174 (RW)
0x1de: frame_vm_group_bin_13711 (RW)
0x1df: frame_vm_group_bin_16218 (RW)
0x1e0: frame_vm_group_bin_9028 (RW)
0x1e1: frame_vm_group_bin_1840 (RW)
0x1e2: frame_vm_group_bin_17941 (RW)
0x1e3: frame_vm_group_bin_10848 (RW)
0x1e4: frame_vm_group_bin_3663 (RW)
0x1e5: frame_vm_group_bin_19763 (RW)
0x1e6: frame_vm_group_bin_12591 (RW)
0x1e7: frame_vm_group_bin_5499 (RW)
0x1e8: frame_vm_group_bin_21596 (RW)
0x1e9: frame_vm_group_bin_14420 (RW)
0x1e: frame_vm_group_bin_18616 (RW)
0x1ea: frame_vm_group_bin_7207 (RW)
0x1eb: frame_vm_group_bin_18357 (RW)
0x1ec: frame_vm_group_bin_16244 (RW)
0x1ed: frame_vm_group_bin_9061 (RW)
0x1ee: frame_vm_group_bin_1873 (RW)
0x1ef: frame_vm_group_bin_17973 (RW)
0x1f0: frame_vm_group_bin_10880 (RW)
0x1f1: frame_vm_group_bin_3696 (RW)
0x1f2: frame_vm_group_bin_19796 (RW)
0x1f3: frame_vm_group_bin_12624 (RW)
0x1f4: frame_vm_group_bin_5531 (RW)
0x1f5: frame_vm_group_bin_21629 (RW)
0x1f6: frame_vm_group_bin_14453 (RW)
0x1f7: frame_vm_group_bin_7240 (RW)
0x1f8: frame_vm_group_bin_23095 (RW)
0x1f9: frame_vm_group_bin_16271 (RW)
0x1f: frame_vm_group_bin_11552 (RW)
0x1fa: frame_vm_group_bin_9095 (RW)
0x1fb: frame_vm_group_bin_1907 (RW)
0x1fc: frame_vm_group_bin_18005 (RW)
0x1fd: frame_vm_group_bin_10915 (RW)
0x1fe: frame_vm_group_bin_3730 (RW)
0x1ff: frame_vm_group_bin_19830 (RW)
0x20: frame_vm_group_bin_4370 (RW)
0x21: frame_vm_group_bin_20466 (RW)
0x22: frame_vm_group_bin_13269 (RW)
0x23: frame_vm_group_bin_6096 (RW)
0x24: frame_vm_group_bin_22276 (RW)
0x25: frame_vm_group_bin_15105 (RW)
0x26: frame_vm_group_bin_7911 (RW)
0x27: frame_vm_group_bin_0747 (RW)
0x28: frame_vm_group_bin_16941 (RW)
0x29: frame_vm_group_bin_9733 (RW)
0x2: frame_vm_group_bin_9634 (RW)
0x2a: frame_vm_group_bin_2572 (RW)
0x2b: frame_vm_group_bin_18648 (RW)
0x2c: frame_vm_group_bin_11580 (RW)
0x2d: frame_vm_group_bin_4403 (RW)
0x2e: frame_vm_group_bin_20499 (RW)
0x2f: frame_vm_group_bin_13302 (RW)
0x30: frame_vm_group_bin_6127 (RW)
0x31: frame_vm_group_bin_22309 (RW)
0x32: frame_vm_group_bin_15131 (RW)
0x33: frame_vm_group_bin_7945 (RW)
0x34: frame_vm_group_bin_0780 (RW)
0x35: frame_vm_group_bin_16974 (RW)
0x36: frame_vm_group_bin_9766 (RW)
0x37: frame_vm_group_bin_2605 (RW)
0x38: frame_vm_group_bin_18681 (RW)
0x39: frame_vm_group_bin_11604 (RW)
0x3: frame_vm_group_bin_2472 (RW)
0x3a: frame_vm_group_bin_4437 (RW)
0x3b: frame_vm_group_bin_20533 (RW)
0x3c: frame_vm_group_bin_13335 (RW)
0x3d: frame_vm_group_bin_6160 (RW)
0x3e: frame_vm_group_bin_22342 (RW)
0x3f: frame_vm_group_bin_15158 (RW)
0x40: frame_vm_group_bin_7979 (RW)
0x41: frame_vm_group_bin_0813 (RW)
0x42: frame_vm_group_bin_17008 (RW)
0x43: frame_vm_group_bin_9800 (RW)
0x44: frame_vm_group_bin_2639 (RW)
0x45: frame_vm_group_bin_18714 (RW)
0x46: frame_vm_group_bin_4340 (RW)
0x47: frame_vm_group_bin_4470 (RW)
0x48: frame_vm_group_bin_20566 (RW)
0x49: frame_vm_group_bin_13368 (RW)
0x4: frame_vm_group_bin_18553 (RW)
0x4a: frame_vm_group_bin_6192 (RW)
0x4b: frame_vm_group_bin_22375 (RW)
0x4c: frame_vm_group_bin_15191 (RW)
0x4d: frame_vm_group_bin_8009 (RW)
0x4e: frame_vm_group_bin_0846 (RW)
0x4f: frame_vm_group_bin_17041 (RW)
0x50: frame_vm_group_bin_9833 (RW)
0x51: frame_vm_group_bin_2672 (RW)
0x52: frame_vm_group_bin_18745 (RW)
0x53: frame_vm_group_bin_20769 (RW)
0x54: frame_vm_group_bin_4503 (RW)
0x55: frame_vm_group_bin_20599 (RW)
0x56: frame_vm_group_bin_13399 (RW)
0x57: frame_vm_group_bin_15044 (RW)
0x58: frame_vm_group_bin_22408 (RW)
0x59: frame_vm_group_bin_15225 (RW)
0x5: frame_vm_group_bin_11485 (RW)
0x5a: frame_vm_group_bin_8038 (RW)
0x5b: frame_vm_group_bin_0880 (RW)
0x5c: frame_vm_group_bin_17075 (RW)
0x5d: frame_vm_group_bin_9867 (RW)
0x5e: frame_vm_group_bin_2706 (RW)
0x5f: frame_vm_group_bin_18779 (RW)
0x60: frame_vm_group_bin_11675 (RW)
0x61: frame_vm_group_bin_4537 (RW)
0x62: frame_vm_group_bin_20633 (RW)
0x63: frame_vm_group_bin_13433 (RW)
0x64: frame_vm_group_bin_6249 (RW)
0x65: frame_vm_group_bin_22441 (RW)
0x66: frame_vm_group_bin_15259 (RW)
0x67: frame_vm_group_bin_8069 (RW)
0x68: frame_vm_group_bin_0913 (RW)
0x69: frame_vm_group_bin_17108 (RW)
0x6: frame_vm_group_bin_4301 (RW)
0x6a: frame_vm_group_bin_9899 (RW)
0x6b: frame_vm_group_bin_2739 (RW)
0x6c: frame_vm_group_bin_18812 (RW)
0x6d: frame_vm_group_bin_11702 (RW)
0x6e: frame_vm_group_bin_4568 (RW)
0x6f: frame_vm_group_bin_20665 (RW)
0x70: frame_vm_group_bin_13466 (RW)
0x71: frame_vm_group_bin_6281 (RW)
0x72: frame_vm_group_bin_22474 (RW)
0x73: frame_vm_group_bin_15291 (RW)
0x74: frame_vm_group_bin_8101 (RW)
0x75: frame_vm_group_bin_0946 (RW)
0x76: frame_vm_group_bin_17141 (RW)
0x77: frame_vm_group_bin_9932 (RW)
0x78: frame_vm_group_bin_2772 (RW)
0x79: frame_vm_group_bin_18846 (RW)
0x7: frame_vm_group_bin_20399 (RW)
0x7a: frame_vm_group_bin_11501 (RW)
0x7b: frame_vm_group_bin_4592 (RW)
0x7c: frame_vm_group_bin_20699 (RW)
0x7d: frame_vm_group_bin_13500 (RW)
0x7e: frame_vm_group_bin_6315 (RW)
0x7f: frame_vm_group_bin_22508 (RW)
0x80: frame_vm_group_bin_15325 (RW)
0x81: frame_vm_group_bin_8134 (RW)
0x82: frame_vm_group_bin_0980 (RW)
0x83: frame_vm_group_bin_17173 (RW)
0x84: frame_vm_group_bin_9964 (RW)
0x85: frame_vm_group_bin_2806 (RW)
0x86: frame_vm_group_bin_18880 (RW)
0x87: frame_vm_group_bin_16145 (RW)
0x88: frame_vm_group_bin_4616 (RW)
0x89: frame_vm_group_bin_20732 (RW)
0x8: frame_vm_group_bin_13202 (RW)
0x8a: frame_vm_group_bin_13533 (RW)
0x8b: frame_vm_group_bin_6347 (RW)
0x8c: frame_vm_group_bin_22540 (RW)
0x8d: frame_vm_group_bin_15358 (RW)
0x8e: frame_vm_group_bin_8167 (RW)
0x8f: frame_vm_group_bin_1012 (RW)
0x90: frame_vm_group_bin_17204 (RW)
0x91: frame_vm_group_bin_9997 (RW)
0x92: frame_vm_group_bin_2839 (RW)
0x93: frame_vm_group_bin_18913 (RW)
0x94: frame_vm_group_bin_20792 (RW)
0x95: frame_vm_group_bin_4644 (RW)
0x96: frame_vm_group_bin_20765 (RW)
0x97: frame_vm_group_bin_13566 (RW)
0x98: frame_vm_group_bin_6379 (RW)
0x99: frame_vm_group_bin_22573 (RW)
0x9: frame_vm_group_bin_10363 (RW)
0x9a: frame_vm_group_bin_15392 (RW)
0x9b: frame_vm_group_bin_8201 (RW)
0x9c: frame_vm_group_bin_1037 (RW)
0x9d: frame_vm_group_bin_17237 (RW)
0x9e: frame_vm_group_bin_10031 (RW)
0x9f: frame_vm_group_bin_2874 (RW)
0xa0: frame_vm_group_bin_18946 (RW)
0xa1: frame_vm_group_bin_11803 (RW)
0xa2: frame_vm_group_bin_4677 (RW)
0xa3: frame_vm_group_bin_20799 (RW)
0xa4: frame_vm_group_bin_13600 (RW)
0xa5: frame_vm_group_bin_6410 (RW)
0xa6: frame_vm_group_bin_22607 (RW)
0xa7: frame_vm_group_bin_15425 (RW)
0xa8: frame_vm_group_bin_8234 (RW)
0xa9: frame_vm_group_bin_1058 (RW)
0xa: frame_vm_group_bin_22210 (RW)
0xaa: frame_vm_group_bin_17270 (RW)
0xab: frame_vm_group_bin_10064 (RW)
0xac: frame_vm_group_bin_2907 (RW)
0xad: frame_vm_group_bin_18977 (RW)
0xae: frame_vm_group_bin_6781 (RW)
0xaf: frame_vm_group_bin_4709 (RW)
0xb0: frame_vm_group_bin_20831 (RW)
0xb1: frame_vm_group_bin_13633 (RW)
0xb2: frame_vm_group_bin_6443 (RW)
0xb3: frame_vm_group_bin_22640 (RW)
0xb4: frame_vm_group_bin_15458 (RW)
0xb5: frame_vm_group_bin_8267 (RW)
0xb6: frame_vm_group_bin_1082 (RW)
0xb7: frame_vm_group_bin_17303 (RW)
0xb8: frame_vm_group_bin_10097 (RW)
0xb9: frame_vm_group_bin_2940 (RW)
0xb: frame_vm_group_bin_15053 (RW)
0xba: frame_vm_group_bin_19011 (RW)
0xbb: frame_vm_group_bin_11865 (RW)
0xbc: frame_vm_group_bin_4742 (RW)
0xbd: frame_vm_group_bin_20860 (RW)
0xbe: frame_vm_group_bin_13666 (RW)
0xbf: frame_vm_group_bin_6477 (RW)
0xc0: frame_vm_group_bin_22674 (RW)
0xc1: frame_vm_group_bin_15492 (RW)
0xc2: frame_vm_group_bin_8300 (RW)
0xc3: frame_vm_group_bin_1112 (RW)
0xc4: frame_vm_group_bin_17337 (RW)
0xc5: frame_vm_group_bin_10131 (RW)
0xc6: frame_vm_group_bin_2974 (RW)
0xc7: frame_vm_group_bin_19044 (RW)
0xc8: frame_vm_group_bin_16170 (RW)
0xc9: frame_vm_group_bin_4775 (RW)
0xc: frame_vm_group_bin_7844 (RW)
0xca: frame_vm_group_bin_20884 (RW)
0xcb: frame_vm_group_bin_13699 (RW)
0xcc: frame_vm_group_bin_6510 (RW)
0xcd: frame_vm_group_bin_22707 (RW)
0xce: frame_vm_group_bin_15524 (RW)
0xcf: frame_vm_group_bin_8333 (RW)
0xd0: frame_vm_group_bin_1144 (RW)
0xd1: frame_vm_group_bin_17369 (RW)
0xd2: frame_vm_group_bin_10166 (RW)
0xd3: frame_vm_group_bin_3007 (RW)
0xd4: frame_vm_group_bin_19077 (RW)
0xd5: frame_vm_group_bin_11916 (RW)
0xd6: frame_vm_group_bin_4808 (RW)
0xd7: frame_vm_group_bin_20912 (RW)
0xd8: frame_vm_group_bin_13731 (RW)
0xd9: frame_vm_group_bin_6543 (RW)
0xd: frame_vm_group_bin_0680 (RW)
0xda: frame_vm_group_bin_22741 (RW)
0xdb: frame_vm_group_bin_15557 (RW)
0xdc: frame_vm_group_bin_8367 (RW)
0xdd: frame_vm_group_bin_1178 (RW)
0xde: frame_vm_group_bin_17400 (RW)
0xdf: frame_vm_group_bin_10200 (RW)
0xe0: frame_vm_group_bin_3041 (RW)
0xe1: frame_vm_group_bin_19110 (RW)
0xe2: frame_vm_group_bin_11946 (RW)
0xe3: frame_vm_group_bin_4841 (RW)
0xe4: frame_vm_group_bin_20942 (RW)
0xe5: frame_vm_group_bin_13766 (RW)
0xe6: frame_vm_group_bin_6577 (RW)
0xe7: frame_vm_group_bin_22773 (RW)
0xe8: frame_vm_group_bin_15590 (RW)
0xe9: frame_vm_group_bin_8400 (RW)
0xe: frame_vm_group_bin_16875 (RW)
0xea: frame_vm_group_bin_1211 (RW)
0xeb: frame_vm_group_bin_17425 (RW)
0xec: frame_vm_group_bin_10233 (RW)
0xed: frame_vm_group_bin_3074 (RW)
0xee: frame_vm_group_bin_19142 (RW)
0xef: frame_vm_group_bin_11979 (RW)
0xf0: frame_vm_group_bin_4874 (RW)
0xf1: frame_vm_group_bin_20967 (RW)
0xf2: frame_vm_group_bin_13799 (RW)
0xf3: frame_vm_group_bin_6610 (RW)
0xf4: frame_vm_group_bin_22806 (RW)
0xf5: frame_vm_group_bin_15623 (RW)
0xf6: frame_vm_group_bin_8433 (RW)
0xf7: frame_vm_group_bin_1244 (RW)
0xf8: frame_vm_group_bin_17450 (RW)
0xf9: frame_vm_group_bin_10266 (RW)
0xf: frame_vm_group_bin_9667 (RW)
0xfa: frame_vm_group_bin_3108 (RW)
0xfb: frame_vm_group_bin_19176 (RW)
0xfc: frame_vm_group_bin_12012 (RW)
0xfd: frame_vm_group_bin_4908 (RW)
0xfe: frame_vm_group_bin_21001 (RW)
0xff: frame_vm_group_bin_13831 (RW)
}
pt_vm_group_bin_0031 {
0x0: frame_vm_group_bin_18476 (RW)
0x100: frame_vm_group_bin_1181 (RW)
0x101: frame_vm_group_bin_17403 (RW)
0x102: frame_vm_group_bin_10203 (RW)
0x103: frame_vm_group_bin_3044 (RW)
0x104: frame_vm_group_bin_19113 (RW)
0x105: frame_vm_group_bin_11949 (RW)
0x106: frame_vm_group_bin_4844 (RW)
0x107: frame_vm_group_bin_7338 (RW)
0x108: frame_vm_group_bin_13769 (RW)
0x109: frame_vm_group_bin_6580 (RW)
0x10: frame_vm_group_bin_20335 (RW)
0x10a: frame_vm_group_bin_22776 (RW)
0x10b: frame_vm_group_bin_15593 (RW)
0x10c: frame_vm_group_bin_8403 (RW)
0x10d: frame_vm_group_bin_1214 (RW)
0x10e: frame_vm_group_bin_20650 (RW)
0x10f: frame_vm_group_bin_10236 (RW)
0x110: frame_vm_group_bin_3077 (RW)
0x111: frame_vm_group_bin_19145 (RW)
0x112: frame_vm_group_bin_11982 (RW)
0x113: frame_vm_group_bin_4877 (RW)
0x114: frame_vm_group_bin_20970 (RW)
0x115: frame_vm_group_bin_13802 (RW)
0x116: frame_vm_group_bin_6613 (RW)
0x117: frame_vm_group_bin_22809 (RW)
0x118: frame_vm_group_bin_15626 (RW)
0x119: frame_vm_group_bin_8436 (RW)
0x11: frame_vm_group_bin_13138 (RW)
0x11a: frame_vm_group_bin_1248 (RW)
0x11b: frame_vm_group_bin_19574 (RW)
0x11c: frame_vm_group_bin_10270 (RW)
0x11d: frame_vm_group_bin_3111 (RW)
0x11e: frame_vm_group_bin_19179 (RW)
0x11f: frame_vm_group_bin_12014 (RW)
0x120: frame_vm_group_bin_4911 (RW)
0x121: frame_vm_group_bin_21004 (RW)
0x122: frame_vm_group_bin_13834 (RW)
0x123: frame_vm_group_bin_6647 (RW)
0x124: frame_vm_group_bin_22843 (RW)
0x125: frame_vm_group_bin_15660 (RW)
0x126: frame_vm_group_bin_8470 (RW)
0x127: frame_vm_group_bin_1278 (RW)
0x128: frame_vm_group_bin_6640 (RW)
0x129: frame_vm_group_bin_10303 (RW)
0x12: frame_vm_group_bin_5985 (RW)
0x12a: frame_vm_group_bin_3143 (RW)
0x12b: frame_vm_group_bin_19212 (RW)
0x12c: frame_vm_group_bin_12044 (RW)
0x12d: frame_vm_group_bin_4942 (RW)
0x12e: frame_vm_group_bin_21037 (RW)
0x12f: frame_vm_group_bin_19919 (RW)
0x130: frame_vm_group_bin_6680 (RW)
0x131: frame_vm_group_bin_22876 (RW)
0x132: frame_vm_group_bin_15693 (RW)
0x133: frame_vm_group_bin_8503 (RW)
0x134: frame_vm_group_bin_1311 (RW)
0x135: frame_vm_group_bin_17494 (RW)
0x136: frame_vm_group_bin_10336 (RW)
0x137: frame_vm_group_bin_3176 (RW)
0x138: frame_vm_group_bin_19245 (RW)
0x139: frame_vm_group_bin_12072 (RW)
0x13: frame_vm_group_bin_22146 (RW)
0x13a: frame_vm_group_bin_4974 (RW)
0x13b: frame_vm_group_bin_21072 (RW)
0x13c: frame_vm_group_bin_13894 (RW)
0x13d: frame_vm_group_bin_23208 (RW)
0x13e: frame_vm_group_bin_22910 (RW)
0x13f: frame_vm_group_bin_15727 (RW)
0x140: frame_vm_group_bin_8536 (RW)
0x141: frame_vm_group_bin_1344 (RW)
0x142: frame_vm_group_bin_17520 (RW)
0x143: frame_vm_group_bin_10370 (RW)
0x144: frame_vm_group_bin_3210 (RW)
0x145: frame_vm_group_bin_19279 (RW)
0x146: frame_vm_group_bin_12106 (RW)
0x147: frame_vm_group_bin_5007 (RW)
0x148: frame_vm_group_bin_21105 (RW)
0x149: frame_vm_group_bin_13927 (RW)
0x14: frame_vm_group_bin_14997 (RW)
0x14a: frame_vm_group_bin_6746 (RW)
0x14b: frame_vm_group_bin_22943 (RW)
0x14c: frame_vm_group_bin_15760 (RW)
0x14d: frame_vm_group_bin_8567 (RW)
0x14e: frame_vm_group_bin_1378 (RW)
0x14f: frame_vm_group_bin_17545 (RW)
0x150: frame_vm_group_bin_10399 (RW)
0x151: frame_vm_group_bin_3242 (RW)
0x152: frame_vm_group_bin_19312 (RW)
0x153: frame_vm_group_bin_12138 (RW)
0x154: frame_vm_group_bin_5040 (RW)
0x155: frame_vm_group_bin_21138 (RW)
0x156: frame_vm_group_bin_13960 (RW)
0x157: frame_vm_group_bin_6778 (RW)
0x158: frame_vm_group_bin_22975 (RW)
0x159: frame_vm_group_bin_15793 (RW)
0x15: frame_vm_group_bin_7781 (RW)
0x15a: frame_vm_group_bin_4929 (RW)
0x15b: frame_vm_group_bin_1412 (RW)
0x15c: frame_vm_group_bin_17568 (RW)
0x15d: frame_vm_group_bin_10426 (RW)
0x15e: frame_vm_group_bin_3276 (RW)
0x15f: frame_vm_group_bin_19346 (RW)
0x160: frame_vm_group_bin_12169 (RW)
0x161: frame_vm_group_bin_5075 (RW)
0x162: frame_vm_group_bin_21171 (RW)
0x163: frame_vm_group_bin_13994 (RW)
0x164: frame_vm_group_bin_6811 (RW)
0x165: frame_vm_group_bin_23008 (RW)
0x166: frame_vm_group_bin_15825 (RW)
0x167: frame_vm_group_bin_8633 (RW)
0x168: frame_vm_group_bin_1445 (RW)
0x169: frame_vm_group_bin_17591 (RW)
0x16: frame_vm_group_bin_0617 (RW)
0x16a: frame_vm_group_bin_10456 (RW)
0x16b: frame_vm_group_bin_3309 (RW)
0x16c: frame_vm_group_bin_19379 (RW)
0x16d: frame_vm_group_bin_12201 (RW)
0x16e: frame_vm_group_bin_5108 (RW)
0x16f: frame_vm_group_bin_21204 (RW)
0x170: frame_vm_group_bin_14027 (RW)
0x171: frame_vm_group_bin_6840 (RW)
0x172: frame_vm_group_bin_23041 (RW)
0x173: frame_vm_group_bin_15858 (RW)
0x174: frame_vm_group_bin_8666 (RW)
0x175: frame_vm_group_bin_1478 (RW)
0x176: frame_vm_group_bin_17618 (RW)
0x177: frame_vm_group_bin_10489 (RW)
0x178: frame_vm_group_bin_3342 (RW)
0x179: frame_vm_group_bin_19412 (RW)
0x17: frame_vm_group_bin_16812 (RW)
0x17a: frame_vm_group_bin_12231 (RW)
0x17b: frame_vm_group_bin_5142 (RW)
0x17c: frame_vm_group_bin_21238 (RW)
0x17d: frame_vm_group_bin_14061 (RW)
0x17e: frame_vm_group_bin_6868 (RW)
0x17f: frame_vm_group_bin_23075 (RW)
0x180: frame_vm_group_bin_15892 (RW)
0x181: frame_vm_group_bin_8701 (RW)
0x182: frame_vm_group_bin_1512 (RW)
0x183: frame_vm_group_bin_17652 (RW)
0x184: frame_vm_group_bin_10522 (RW)
0x185: frame_vm_group_bin_3375 (RW)
0x186: frame_vm_group_bin_19443 (RW)
0x187: frame_vm_group_bin_12264 (RW)
0x188: frame_vm_group_bin_5175 (RW)
0x189: frame_vm_group_bin_21271 (RW)
0x18: frame_vm_group_bin_9603 (RW)
0x18a: frame_vm_group_bin_14094 (RW)
0x18b: frame_vm_group_bin_4591 (RW)
0x18c: frame_vm_group_bin_23108 (RW)
0x18d: frame_vm_group_bin_15925 (RW)
0x18e: frame_vm_group_bin_8734 (RW)
0x18f: frame_vm_group_bin_1545 (RW)
0x190: frame_vm_group_bin_17683 (RW)
0x191: frame_vm_group_bin_10555 (RW)
0x192: frame_vm_group_bin_3404 (RW)
0x193: frame_vm_group_bin_19475 (RW)
0x194: frame_vm_group_bin_12297 (RW)
0x195: frame_vm_group_bin_5208 (RW)
0x196: frame_vm_group_bin_21304 (RW)
0x197: frame_vm_group_bin_14127 (RW)
0x198: frame_vm_group_bin_6917 (RW)
0x199: frame_vm_group_bin_7761 (RW)
0x19: frame_vm_group_bin_2442 (RW)
0x19a: frame_vm_group_bin_15959 (RW)
0x19b: frame_vm_group_bin_8768 (RW)
0x19c: frame_vm_group_bin_1579 (RW)
0x19d: frame_vm_group_bin_17711 (RW)
0x19e: frame_vm_group_bin_10589 (RW)
0x19f: frame_vm_group_bin_3429 (RW)
0x1: frame_vm_group_bin_11389 (RW)
0x1a0: frame_vm_group_bin_19509 (RW)
0x1a1: frame_vm_group_bin_12330 (RW)
0x1a2: frame_vm_group_bin_5242 (RW)
0x1a3: frame_vm_group_bin_21336 (RW)
0x1a4: frame_vm_group_bin_14161 (RW)
0x1a5: frame_vm_group_bin_6948 (RW)
0x1a6: frame_vm_group_bin_23174 (RW)
0x1a7: frame_vm_group_bin_15994 (RW)
0x1a8: frame_vm_group_bin_8801 (RW)
0x1a9: frame_vm_group_bin_1612 (RW)
0x1a: frame_vm_group_bin_18529 (RW)
0x1aa: frame_vm_group_bin_17737 (RW)
0x1ab: frame_vm_group_bin_10622 (RW)
0x1ac: frame_vm_group_bin_3870 (RW)
0x1ad: frame_vm_group_bin_19542 (RW)
0x1ae: frame_vm_group_bin_12363 (RW)
0x1af: frame_vm_group_bin_5275 (RW)
0x1b0: frame_vm_group_bin_21369 (RW)
0x1b1: frame_vm_group_bin_14193 (RW)
0x1b2: frame_vm_group_bin_6980 (RW)
0x1b3: frame_vm_group_bin_23205 (RW)
0x1b4: frame_vm_group_bin_16027 (RW)
0x1b5: frame_vm_group_bin_8834 (RW)
0x1b6: frame_vm_group_bin_1645 (RW)
0x1b7: frame_vm_group_bin_17765 (RW)
0x1b8: frame_vm_group_bin_10654 (RW)
0x1b9: frame_vm_group_bin_3477 (RW)
0x1b: frame_vm_group_bin_11455 (RW)
0x1ba: frame_vm_group_bin_19577 (RW)
0x1bb: frame_vm_group_bin_12397 (RW)
0x1bc: frame_vm_group_bin_5309 (RW)
0x1bd: frame_vm_group_bin_21403 (RW)
0x1be: frame_vm_group_bin_14227 (RW)
0x1bf: frame_vm_group_bin_7014 (RW)
0x1c0: frame_vm_group_bin_21800 (RW)
0x1c1: frame_vm_group_bin_16061 (RW)
0x1c2: frame_vm_group_bin_8867 (RW)
0x1c3: frame_vm_group_bin_1679 (RW)
0x1c4: frame_vm_group_bin_17796 (RW)
0x1c5: frame_vm_group_bin_10687 (RW)
0x1c6: frame_vm_group_bin_3505 (RW)
0x1c7: frame_vm_group_bin_19610 (RW)
0x1c8: frame_vm_group_bin_12430 (RW)
0x1c9: frame_vm_group_bin_5340 (RW)
0x1c: frame_vm_group_bin_4271 (RW)
0x1ca: frame_vm_group_bin_21435 (RW)
0x1cb: frame_vm_group_bin_14259 (RW)
0x1cc: frame_vm_group_bin_7046 (RW)
0x1cd: frame_vm_group_bin_3179 (RW)
0x1ce: frame_vm_group_bin_16093 (RW)
0x1cf: frame_vm_group_bin_8899 (RW)
0x1d0: frame_vm_group_bin_1711 (RW)
0x1d1: frame_vm_group_bin_17826 (RW)
0x1d2: frame_vm_group_bin_10719 (RW)
0x1d3: frame_vm_group_bin_3533 (RW)
0x1d4: frame_vm_group_bin_19641 (RW)
0x1d5: frame_vm_group_bin_12461 (RW)
0x1d6: frame_vm_group_bin_5371 (RW)
0x1d7: frame_vm_group_bin_21467 (RW)
0x1d8: frame_vm_group_bin_10701 (RW)
0x1d9: frame_vm_group_bin_7077 (RW)
0x1d: frame_vm_group_bin_20369 (RW)
0x1da: frame_vm_group_bin_0016 (RW)
0x1db: frame_vm_group_bin_16126 (RW)
0x1dc: frame_vm_group_bin_8932 (RW)
0x1dd: frame_vm_group_bin_1744 (RW)
0x1de: frame_vm_group_bin_17854 (RW)
0x1df: frame_vm_group_bin_10752 (RW)
0x1e0: frame_vm_group_bin_3565 (RW)
0x1e1: frame_vm_group_bin_19669 (RW)
0x1e2: frame_vm_group_bin_12494 (RW)
0x1e3: frame_vm_group_bin_5404 (RW)
0x1e4: frame_vm_group_bin_21499 (RW)
0x1e5: frame_vm_group_bin_14323 (RW)
0x1e6: frame_vm_group_bin_7109 (RW)
0x1e7: frame_vm_group_bin_12442 (RW)
0x1e8: frame_vm_group_bin_16157 (RW)
0x1e9: frame_vm_group_bin_8964 (RW)
0x1e: frame_vm_group_bin_13172 (RW)
0x1ea: frame_vm_group_bin_1776 (RW)
0x1eb: frame_vm_group_bin_17880 (RW)
0x1ec: frame_vm_group_bin_10784 (RW)
0x1ed: frame_vm_group_bin_3599 (RW)
0x1ee: frame_vm_group_bin_19699 (RW)
0x1ef: frame_vm_group_bin_12527 (RW)
0x1f0: frame_vm_group_bin_5437 (RW)
0x1f1: frame_vm_group_bin_21532 (RW)
0x1f2: frame_vm_group_bin_14356 (RW)
0x1f3: frame_vm_group_bin_7141 (RW)
0x1f4: frame_vm_group_bin_0059 (RW)
0x1f5: frame_vm_group_bin_16190 (RW)
0x1f6: frame_vm_group_bin_8997 (RW)
0x1f7: frame_vm_group_bin_1809 (RW)
0x1f8: frame_vm_group_bin_17911 (RW)
0x1f9: frame_vm_group_bin_10817 (RW)
0x1f: frame_vm_group_bin_6016 (RW)
0x1fa: frame_vm_group_bin_3633 (RW)
0x1fb: frame_vm_group_bin_19733 (RW)
0x1fc: frame_vm_group_bin_12561 (RW)
0x1fd: frame_vm_group_bin_5470 (RW)
0x1fe: frame_vm_group_bin_21566 (RW)
0x1ff: frame_vm_group_bin_14390 (RW)
0x20: frame_vm_group_bin_22180 (RW)
0x21: frame_vm_group_bin_15031 (RW)
0x22: frame_vm_group_bin_7815 (RW)
0x23: frame_vm_group_bin_0650 (RW)
0x24: frame_vm_group_bin_16846 (RW)
0x25: frame_vm_group_bin_9637 (RW)
0x26: frame_vm_group_bin_2475 (RW)
0x27: frame_vm_group_bin_2278 (RW)
0x28: frame_vm_group_bin_11488 (RW)
0x29: frame_vm_group_bin_4304 (RW)
0x2: frame_vm_group_bin_4204 (RW)
0x2a: frame_vm_group_bin_20402 (RW)
0x2b: frame_vm_group_bin_13205 (RW)
0x2c: frame_vm_group_bin_6044 (RW)
0x2d: frame_vm_group_bin_22213 (RW)
0x2e: frame_vm_group_bin_15056 (RW)
0x2f: frame_vm_group_bin_7847 (RW)
0x30: frame_vm_group_bin_0683 (RW)
0x31: frame_vm_group_bin_16878 (RW)
0x32: frame_vm_group_bin_9670 (RW)
0x33: frame_vm_group_bin_2508 (RW)
0x34: frame_vm_group_bin_18585 (RW)
0x35: frame_vm_group_bin_11521 (RW)
0x36: frame_vm_group_bin_4337 (RW)
0x37: frame_vm_group_bin_20435 (RW)
0x38: frame_vm_group_bin_13238 (RW)
0x39: frame_vm_group_bin_6068 (RW)
0x3: frame_vm_group_bin_20300 (RW)
0x3a: frame_vm_group_bin_22247 (RW)
0x3b: frame_vm_group_bin_15081 (RW)
0x3c: frame_vm_group_bin_7881 (RW)
0x3d: frame_vm_group_bin_0717 (RW)
0x3e: frame_vm_group_bin_16911 (RW)
0x3f: frame_vm_group_bin_9703 (RW)
0x40: frame_vm_group_bin_2542 (RW)
0x41: frame_vm_group_bin_18619 (RW)
0x42: frame_vm_group_bin_11555 (RW)
0x43: frame_vm_group_bin_4373 (RW)
0x44: frame_vm_group_bin_20469 (RW)
0x45: frame_vm_group_bin_13272 (RW)
0x46: frame_vm_group_bin_6099 (RW)
0x47: frame_vm_group_bin_22279 (RW)
0x48: frame_vm_group_bin_1553 (RW)
0x49: frame_vm_group_bin_7914 (RW)
0x4: frame_vm_group_bin_13105 (RW)
0x4a: frame_vm_group_bin_0750 (RW)
0x4b: frame_vm_group_bin_16944 (RW)
0x4c: frame_vm_group_bin_9736 (RW)
0x4d: frame_vm_group_bin_2575 (RW)
0x4e: frame_vm_group_bin_18651 (RW)
0x4f: frame_vm_group_bin_11583 (RW)
0x50: frame_vm_group_bin_4406 (RW)
0x51: frame_vm_group_bin_20502 (RW)
0x52: frame_vm_group_bin_13305 (RW)
0x53: frame_vm_group_bin_6130 (RW)
0x54: frame_vm_group_bin_22312 (RW)
0x55: frame_vm_group_bin_6204 (RW)
0x56: frame_vm_group_bin_7948 (RW)
0x57: frame_vm_group_bin_0783 (RW)
0x58: frame_vm_group_bin_16977 (RW)
0x59: frame_vm_group_bin_9769 (RW)
0x5: frame_vm_group_bin_5956 (RW)
0x5a: frame_vm_group_bin_2609 (RW)
0x5b: frame_vm_group_bin_18685 (RW)
0x5c: frame_vm_group_bin_11608 (RW)
0x5d: frame_vm_group_bin_4440 (RW)
0x5e: frame_vm_group_bin_20536 (RW)
0x5f: frame_vm_group_bin_13338 (RW)
0x60: frame_vm_group_bin_6163 (RW)
0x61: frame_vm_group_bin_22345 (RW)
0x62: frame_vm_group_bin_15161 (RW)
0x63: frame_vm_group_bin_7982 (RW)
0x64: frame_vm_group_bin_0816 (RW)
0x65: frame_vm_group_bin_17011 (RW)
0x66: frame_vm_group_bin_9803 (RW)
0x67: frame_vm_group_bin_2642 (RW)
0x68: frame_vm_group_bin_18717 (RW)
0x69: frame_vm_group_bin_6450 (RW)
0x6: frame_vm_group_bin_22113 (RW)
0x6a: frame_vm_group_bin_4473 (RW)
0x6b: frame_vm_group_bin_20569 (RW)
0x6c: frame_vm_group_bin_13371 (RW)
0x6d: frame_vm_group_bin_6194 (RW)
0x6e: frame_vm_group_bin_22378 (RW)
0x6f: frame_vm_group_bin_15194 (RW)
0x70: frame_vm_group_bin_8012 (RW)
0x71: frame_vm_group_bin_0849 (RW)
0x72: frame_vm_group_bin_17044 (RW)
0x73: frame_vm_group_bin_9836 (RW)
0x74: frame_vm_group_bin_2675 (RW)
0x75: frame_vm_group_bin_18748 (RW)
0x76: frame_vm_group_bin_5583 (RW)
0x77: frame_vm_group_bin_4506 (RW)
0x78: frame_vm_group_bin_20602 (RW)
0x79: frame_vm_group_bin_13402 (RW)
0x7: frame_vm_group_bin_14964 (RW)
0x7a: frame_vm_group_bin_6222 (RW)
0x7b: frame_vm_group_bin_22412 (RW)
0x7c: frame_vm_group_bin_15229 (RW)
0x7d: frame_vm_group_bin_8041 (RW)
0x7e: frame_vm_group_bin_0883 (RW)
0x7f: frame_vm_group_bin_17078 (RW)
0x80: frame_vm_group_bin_9870 (RW)
0x81: frame_vm_group_bin_2709 (RW)
0x82: frame_vm_group_bin_18782 (RW)
0x83: frame_vm_group_bin_11677 (RW)
0x84: frame_vm_group_bin_4540 (RW)
0x85: frame_vm_group_bin_20636 (RW)
0x86: frame_vm_group_bin_13436 (RW)
0x87: frame_vm_group_bin_6252 (RW)
0x88: frame_vm_group_bin_22444 (RW)
0x89: frame_vm_group_bin_15262 (RW)
0x8: frame_vm_group_bin_7748 (RW)
0x8a: frame_vm_group_bin_8072 (RW)
0x8b: frame_vm_group_bin_0916 (RW)
0x8c: frame_vm_group_bin_17111 (RW)
0x8d: frame_vm_group_bin_9902 (RW)
0x8e: frame_vm_group_bin_2742 (RW)
0x8f: frame_vm_group_bin_18815 (RW)
0x90: frame_vm_group_bin_11704 (RW)
0x91: frame_vm_group_bin_4571 (RW)
0x92: frame_vm_group_bin_20668 (RW)
0x93: frame_vm_group_bin_13469 (RW)
0x94: frame_vm_group_bin_6284 (RW)
0x95: frame_vm_group_bin_22477 (RW)
0x96: frame_vm_group_bin_15294 (RW)
0x97: frame_vm_group_bin_8104 (RW)
0x98: frame_vm_group_bin_0949 (RW)
0x99: frame_vm_group_bin_17144 (RW)
0x9: frame_vm_group_bin_0584 (RW)
0x9a: frame_vm_group_bin_0505 (RW)
0x9b: frame_vm_group_bin_2776 (RW)
0x9c: frame_vm_group_bin_18850 (RW)
0x9d: frame_vm_group_bin_11730 (RW)
0x9e: frame_vm_group_bin_18052 (RW)
0x9f: frame_vm_group_bin_20702 (RW)
0xa0: frame_vm_group_bin_13503 (RW)
0xa1: frame_vm_group_bin_6317 (RW)
0xa2: frame_vm_group_bin_22511 (RW)
0xa3: frame_vm_group_bin_15328 (RW)
0xa4: frame_vm_group_bin_8137 (RW)
0xa5: frame_vm_group_bin_0983 (RW)
0xa6: frame_vm_group_bin_17176 (RW)
0xa7: frame_vm_group_bin_9967 (RW)
0xa8: frame_vm_group_bin_2809 (RW)
0xa9: frame_vm_group_bin_18883 (RW)
0xa: frame_vm_group_bin_16779 (RW)
0xaa: frame_vm_group_bin_0879 (RW)
0xab: frame_vm_group_bin_22789 (RW)
0xac: frame_vm_group_bin_20735 (RW)
0xad: frame_vm_group_bin_13536 (RW)
0xae: frame_vm_group_bin_6350 (RW)
0xaf: frame_vm_group_bin_22543 (RW)
0xb0: frame_vm_group_bin_15361 (RW)
0xb1: frame_vm_group_bin_8170 (RW)
0xb2: frame_vm_group_bin_1015 (RW)
0xb3: frame_vm_group_bin_17207 (RW)
0xb4: frame_vm_group_bin_10000 (RW)
0xb5: frame_vm_group_bin_2842 (RW)
0xb6: frame_vm_group_bin_18916 (RW)
0xb7: frame_vm_group_bin_11776 (RW)
0xb8: frame_vm_group_bin_4647 (RW)
0xb9: frame_vm_group_bin_20768 (RW)
0xb: frame_vm_group_bin_9570 (RW)
0xba: frame_vm_group_bin_13570 (RW)
0xbb: frame_vm_group_bin_23164 (RW)
0xbc: frame_vm_group_bin_22577 (RW)
0xbd: frame_vm_group_bin_15395 (RW)
0xbe: frame_vm_group_bin_8204 (RW)
0xbf: frame_vm_group_bin_1040 (RW)
0xc0: frame_vm_group_bin_17240 (RW)
0xc1: frame_vm_group_bin_10034 (RW)
0xc2: frame_vm_group_bin_2877 (RW)
0xc3: frame_vm_group_bin_18949 (RW)
0xc4: frame_vm_group_bin_11806 (RW)
0xc5: frame_vm_group_bin_4680 (RW)
0xc6: frame_vm_group_bin_20802 (RW)
0xc7: frame_vm_group_bin_13603 (RW)
0xc8: frame_vm_group_bin_6413 (RW)
0xc9: frame_vm_group_bin_22610 (RW)
0xc: frame_vm_group_bin_2410 (RW)
0xca: frame_vm_group_bin_15428 (RW)
0xcb: frame_vm_group_bin_8237 (RW)
0xcc: frame_vm_group_bin_22063 (RW)
0xcd: frame_vm_group_bin_17273 (RW)
0xce: frame_vm_group_bin_10067 (RW)
0xcf: frame_vm_group_bin_2910 (RW)
0xd0: frame_vm_group_bin_18980 (RW)
0xd1: frame_vm_group_bin_11838 (RW)
0xd2: frame_vm_group_bin_4712 (RW)
0xd3: frame_vm_group_bin_20834 (RW)
0xd4: frame_vm_group_bin_13636 (RW)
0xd5: frame_vm_group_bin_6446 (RW)
0xd6: frame_vm_group_bin_22643 (RW)
0xd7: frame_vm_group_bin_15461 (RW)
0xd8: frame_vm_group_bin_4882 (RW)
0xd9: frame_vm_group_bin_1085 (RW)
0xd: frame_vm_group_bin_16272 (RW)
0xda: frame_vm_group_bin_17307 (RW)
0xdb: frame_vm_group_bin_10101 (RW)
0xdc: frame_vm_group_bin_2944 (RW)
0xdd: frame_vm_group_bin_19014 (RW)
0xde: frame_vm_group_bin_11868 (RW)
0xdf: frame_vm_group_bin_4745 (RW)
0xe0: frame_vm_group_bin_20863 (RW)
0xe1: frame_vm_group_bin_13669 (RW)
0xe2: frame_vm_group_bin_6480 (RW)
0xe3: frame_vm_group_bin_22677 (RW)
0xe4: frame_vm_group_bin_15495 (RW)
0xe5: frame_vm_group_bin_8303 (RW)
0xe6: frame_vm_group_bin_8060 (RW)
0xe7: frame_vm_group_bin_17340 (RW)
0xe8: frame_vm_group_bin_10134 (RW)
0xe9: frame_vm_group_bin_2977 (RW)
0xe: frame_vm_group_bin_11421 (RW)
0xea: frame_vm_group_bin_19047 (RW)
0xeb: frame_vm_group_bin_11892 (RW)
0xec: frame_vm_group_bin_4778 (RW)
0xed: frame_vm_group_bin_21352 (RW)
0xee: frame_vm_group_bin_13702 (RW)
0xef: frame_vm_group_bin_6513 (RW)
0xf0: frame_vm_group_bin_22710 (RW)
0xf1: frame_vm_group_bin_15527 (RW)
0xf2: frame_vm_group_bin_8336 (RW)
0xf3: frame_vm_group_bin_1147 (RW)
0xf4: frame_vm_group_bin_17372 (RW)
0xf5: frame_vm_group_bin_10169 (RW)
0xf6: frame_vm_group_bin_3010 (RW)
0xf7: frame_vm_group_bin_19080 (RW)
0xf8: frame_vm_group_bin_11918 (RW)
0xf9: frame_vm_group_bin_4811 (RW)
0xf: frame_vm_group_bin_4237 (RW)
0xfa: frame_vm_group_bin_20916 (RW)
0xfb: frame_vm_group_bin_13735 (RW)
0xfc: frame_vm_group_bin_6547 (RW)
0xfd: frame_vm_group_bin_22744 (RW)
0xfe: frame_vm_group_bin_15560 (RW)
0xff: frame_vm_group_bin_8370 (RW)
}
pt_vm_group_bin_0033 {
0x0: frame_vm_group_bin_20703 (RW)
0x100: frame_vm_group_bin_17453 (RW)
0x101: frame_vm_group_bin_19510 (RW)
0x102: frame_vm_group_bin_12331 (RW)
0x103: frame_vm_group_bin_5243 (RW)
0x104: frame_vm_group_bin_21337 (RW)
0x105: frame_vm_group_bin_14162 (RW)
0x106: frame_vm_group_bin_6949 (RW)
0x107: frame_vm_group_bin_23175 (RW)
0x108: frame_vm_group_bin_15995 (RW)
0x109: frame_vm_group_bin_8802 (RW)
0x10: frame_vm_group_bin_22544 (RW)
0x10a: frame_vm_group_bin_1613 (RW)
0x10b: frame_vm_group_bin_17738 (RW)
0x10c: frame_vm_group_bin_10623 (RW)
0x10d: frame_vm_group_bin_22082 (RW)
0x10e: frame_vm_group_bin_19543 (RW)
0x10f: frame_vm_group_bin_12364 (RW)
0x110: frame_vm_group_bin_5276 (RW)
0x111: frame_vm_group_bin_21370 (RW)
0x112: frame_vm_group_bin_14194 (RW)
0x113: frame_vm_group_bin_6981 (RW)
0x114: frame_vm_group_bin_23206 (RW)
0x115: frame_vm_group_bin_16028 (RW)
0x116: frame_vm_group_bin_8835 (RW)
0x117: frame_vm_group_bin_1646 (RW)
0x118: frame_vm_group_bin_17766 (RW)
0x119: frame_vm_group_bin_10655 (RW)
0x11: frame_vm_group_bin_15362 (RW)
0x11a: frame_vm_group_bin_3479 (RW)
0x11b: frame_vm_group_bin_19578 (RW)
0x11c: frame_vm_group_bin_12398 (RW)
0x11d: frame_vm_group_bin_5310 (RW)
0x11e: frame_vm_group_bin_21404 (RW)
0x11f: frame_vm_group_bin_14228 (RW)
0x120: frame_vm_group_bin_7015 (RW)
0x121: frame_vm_group_bin_16742 (RW)
0x122: frame_vm_group_bin_16062 (RW)
0x123: frame_vm_group_bin_8868 (RW)
0x124: frame_vm_group_bin_1680 (RW)
0x125: frame_vm_group_bin_17797 (RW)
0x126: frame_vm_group_bin_10688 (RW)
0x127: frame_vm_group_bin_8084 (RW)
0x128: frame_vm_group_bin_19611 (RW)
0x129: frame_vm_group_bin_12431 (RW)
0x12: frame_vm_group_bin_8171 (RW)
0x12a: frame_vm_group_bin_5341 (RW)
0x12b: frame_vm_group_bin_21436 (RW)
0x12c: frame_vm_group_bin_14260 (RW)
0x12d: frame_vm_group_bin_7047 (RW)
0x12e: frame_vm_group_bin_21376 (RW)
0x12f: frame_vm_group_bin_16094 (RW)
0x130: frame_vm_group_bin_8900 (RW)
0x131: frame_vm_group_bin_1712 (RW)
0x132: frame_vm_group_bin_17827 (RW)
0x133: frame_vm_group_bin_10720 (RW)
0x134: frame_vm_group_bin_3534 (RW)
0x135: frame_vm_group_bin_19642 (RW)
0x136: frame_vm_group_bin_12462 (RW)
0x137: frame_vm_group_bin_5372 (RW)
0x138: frame_vm_group_bin_21468 (RW)
0x139: frame_vm_group_bin_14291 (RW)
0x13: frame_vm_group_bin_1016 (RW)
0x13a: frame_vm_group_bin_7079 (RW)
0x13b: frame_vm_group_bin_0017 (RW)
0x13c: frame_vm_group_bin_16127 (RW)
0x13d: frame_vm_group_bin_8933 (RW)
0x13e: frame_vm_group_bin_1745 (RW)
0x13f: frame_vm_group_bin_20293 (RW)
0x140: frame_vm_group_bin_10753 (RW)
0x141: frame_vm_group_bin_3566 (RW)
0x142: frame_vm_group_bin_19670 (RW)
0x143: frame_vm_group_bin_12495 (RW)
0x144: frame_vm_group_bin_5405 (RW)
0x145: frame_vm_group_bin_21500 (RW)
0x146: frame_vm_group_bin_14324 (RW)
0x147: frame_vm_group_bin_7110 (RW)
0x148: frame_vm_group_bin_0035 (RW)
0x149: frame_vm_group_bin_16158 (RW)
0x14: frame_vm_group_bin_17208 (RW)
0x14a: frame_vm_group_bin_8965 (RW)
0x14b: frame_vm_group_bin_1777 (RW)
0x14c: frame_vm_group_bin_17881 (RW)
0x14d: frame_vm_group_bin_10785 (RW)
0x14e: frame_vm_group_bin_3600 (RW)
0x14f: frame_vm_group_bin_19700 (RW)
0x150: frame_vm_group_bin_12528 (RW)
0x151: frame_vm_group_bin_5438 (RW)
0x152: frame_vm_group_bin_21533 (RW)
0x153: frame_vm_group_bin_14357 (RW)
0x154: frame_vm_group_bin_7142 (RW)
0x155: frame_vm_group_bin_0060 (RW)
0x156: frame_vm_group_bin_16191 (RW)
0x157: frame_vm_group_bin_8998 (RW)
0x158: frame_vm_group_bin_1810 (RW)
0x159: frame_vm_group_bin_17912 (RW)
0x15: frame_vm_group_bin_10001 (RW)
0x15a: frame_vm_group_bin_10819 (RW)
0x15b: frame_vm_group_bin_3634 (RW)
0x15c: frame_vm_group_bin_19734 (RW)
0x15d: frame_vm_group_bin_12562 (RW)
0x15e: frame_vm_group_bin_22482 (RW)
0x15f: frame_vm_group_bin_21567 (RW)
0x160: frame_vm_group_bin_14391 (RW)
0x161: frame_vm_group_bin_7178 (RW)
0x162: frame_vm_group_bin_0087 (RW)
0x163: frame_vm_group_bin_15298 (RW)
0x164: frame_vm_group_bin_9032 (RW)
0x165: frame_vm_group_bin_1844 (RW)
0x166: frame_vm_group_bin_17945 (RW)
0x167: frame_vm_group_bin_10852 (RW)
0x168: frame_vm_group_bin_3667 (RW)
0x169: frame_vm_group_bin_19767 (RW)
0x16: frame_vm_group_bin_2843 (RW)
0x16a: frame_vm_group_bin_12595 (RW)
0x16b: frame_vm_group_bin_5503 (RW)
0x16c: frame_vm_group_bin_21600 (RW)
0x16d: frame_vm_group_bin_14424 (RW)
0x16e: frame_vm_group_bin_7211 (RW)
0x16f: frame_vm_group_bin_0112 (RW)
0x170: frame_vm_group_bin_19943 (RW)
0x171: frame_vm_group_bin_9065 (RW)
0x172: frame_vm_group_bin_1877 (RW)
0x173: frame_vm_group_bin_17975 (RW)
0x174: frame_vm_group_bin_10884 (RW)
0x175: frame_vm_group_bin_3700 (RW)
0x176: frame_vm_group_bin_19800 (RW)
0x177: frame_vm_group_bin_12628 (RW)
0x178: frame_vm_group_bin_5535 (RW)
0x179: frame_vm_group_bin_21633 (RW)
0x17: frame_vm_group_bin_18917 (RW)
0x17a: frame_vm_group_bin_14458 (RW)
0x17b: frame_vm_group_bin_7245 (RW)
0x17c: frame_vm_group_bin_0135 (RW)
0x17d: frame_vm_group_bin_16276 (RW)
0x17e: frame_vm_group_bin_9099 (RW)
0x17f: frame_vm_group_bin_1911 (RW)
0x180: frame_vm_group_bin_18009 (RW)
0x181: frame_vm_group_bin_10919 (RW)
0x182: frame_vm_group_bin_3734 (RW)
0x183: frame_vm_group_bin_19834 (RW)
0x184: frame_vm_group_bin_12660 (RW)
0x185: frame_vm_group_bin_5569 (RW)
0x186: frame_vm_group_bin_21667 (RW)
0x187: frame_vm_group_bin_14491 (RW)
0x188: frame_vm_group_bin_7278 (RW)
0x189: frame_vm_group_bin_0156 (RW)
0x18: frame_vm_group_bin_11777 (RW)
0x18a: frame_vm_group_bin_16307 (RW)
0x18b: frame_vm_group_bin_9132 (RW)
0x18c: frame_vm_group_bin_1944 (RW)
0x18d: frame_vm_group_bin_18042 (RW)
0x18e: frame_vm_group_bin_10952 (RW)
0x18f: frame_vm_group_bin_3767 (RW)
0x190: frame_vm_group_bin_19867 (RW)
0x191: frame_vm_group_bin_19224 (RW)
0x192: frame_vm_group_bin_5601 (RW)
0x193: frame_vm_group_bin_21699 (RW)
0x194: frame_vm_group_bin_14525 (RW)
0x195: frame_vm_group_bin_7310 (RW)
0x196: frame_vm_group_bin_0185 (RW)
0x197: frame_vm_group_bin_16339 (RW)
0x198: frame_vm_group_bin_9225 (RW)
0x199: frame_vm_group_bin_1976 (RW)
0x19: frame_vm_group_bin_4648 (RW)
0x19a: frame_vm_group_bin_18075 (RW)
0x19b: frame_vm_group_bin_10985 (RW)
0x19c: frame_vm_group_bin_3800 (RW)
0x19d: frame_vm_group_bin_2047 (RW)
0x19e: frame_vm_group_bin_12709 (RW)
0x19f: frame_vm_group_bin_5633 (RW)
0x1: frame_vm_group_bin_13504 (RW)
0x1a0: frame_vm_group_bin_21733 (RW)
0x1a1: frame_vm_group_bin_14559 (RW)
0x1a2: frame_vm_group_bin_7344 (RW)
0x1a3: frame_vm_group_bin_0217 (RW)
0x1a4: frame_vm_group_bin_16373 (RW)
0x1a5: frame_vm_group_bin_9196 (RW)
0x1a6: frame_vm_group_bin_2010 (RW)
0x1a7: frame_vm_group_bin_18106 (RW)
0x1a8: frame_vm_group_bin_11018 (RW)
0x1a9: frame_vm_group_bin_3833 (RW)
0x1a: frame_vm_group_bin_20770 (RW)
0x1aa: frame_vm_group_bin_19931 (RW)
0x1ab: frame_vm_group_bin_5328 (RW)
0x1ac: frame_vm_group_bin_5666 (RW)
0x1ad: frame_vm_group_bin_21766 (RW)
0x1ae: frame_vm_group_bin_14592 (RW)
0x1af: frame_vm_group_bin_7377 (RW)
0x1b0: frame_vm_group_bin_0242 (RW)
0x1b1: frame_vm_group_bin_16406 (RW)
0x1b2: frame_vm_group_bin_18510 (RW)
0x1b3: frame_vm_group_bin_2043 (RW)
0x1b4: frame_vm_group_bin_18139 (RW)
0x1b5: frame_vm_group_bin_11051 (RW)
0x1b6: frame_vm_group_bin_3866 (RW)
0x1b7: frame_vm_group_bin_19964 (RW)
0x1b8: frame_vm_group_bin_12763 (RW)
0x1b9: frame_vm_group_bin_5699 (RW)
0x1b: frame_vm_group_bin_13571 (RW)
0x1ba: frame_vm_group_bin_7034 (RW)
0x1bb: frame_vm_group_bin_14625 (RW)
0x1bc: frame_vm_group_bin_7411 (RW)
0x1bd: frame_vm_group_bin_0265 (RW)
0x1be: frame_vm_group_bin_16440 (RW)
0x1bf: frame_vm_group_bin_23239 (RW)
0x1c0: frame_vm_group_bin_2077 (RW)
0x1c1: frame_vm_group_bin_18173 (RW)
0x1c2: frame_vm_group_bin_11085 (RW)
0x1c3: frame_vm_group_bin_3900 (RW)
0x1c4: frame_vm_group_bin_19996 (RW)
0x1c5: frame_vm_group_bin_12797 (RW)
0x1c6: frame_vm_group_bin_5733 (RW)
0x1c7: frame_vm_group_bin_21833 (RW)
0x1c8: frame_vm_group_bin_14658 (RW)
0x1c9: frame_vm_group_bin_7444 (RW)
0x1c: frame_vm_group_bin_18004 (RW)
0x1ca: frame_vm_group_bin_0292 (RW)
0x1cb: frame_vm_group_bin_16473 (RW)
0x1cc: frame_vm_group_bin_4609 (RW)
0x1cd: frame_vm_group_bin_2110 (RW)
0x1ce: frame_vm_group_bin_18205 (RW)
0x1cf: frame_vm_group_bin_11118 (RW)
0x1d0: frame_vm_group_bin_3933 (RW)
0x1d1: frame_vm_group_bin_20029 (RW)
0x1d2: frame_vm_group_bin_12829 (RW)
0x1d3: frame_vm_group_bin_17810 (RW)
0x1d4: frame_vm_group_bin_21866 (RW)
0x1d5: frame_vm_group_bin_14691 (RW)
0x1d6: frame_vm_group_bin_7477 (RW)
0x1d7: frame_vm_group_bin_0324 (RW)
0x1d8: frame_vm_group_bin_16506 (RW)
0x1d9: frame_vm_group_bin_9297 (RW)
0x1d: frame_vm_group_bin_22578 (RW)
0x1da: frame_vm_group_bin_2145 (RW)
0x1db: frame_vm_group_bin_18239 (RW)
0x1dc: frame_vm_group_bin_11151 (RW)
0x1dd: frame_vm_group_bin_3966 (RW)
0x1de: frame_vm_group_bin_20063 (RW)
0x1df: frame_vm_group_bin_12863 (RW)
0x1e0: frame_vm_group_bin_22527 (RW)
0x1e1: frame_vm_group_bin_21900 (RW)
0x1e2: frame_vm_group_bin_14725 (RW)
0x1e3: frame_vm_group_bin_7510 (RW)
0x1e4: frame_vm_group_bin_0356 (RW)
0x1e5: frame_vm_group_bin_16540 (RW)
0x1e6: frame_vm_group_bin_9328 (RW)
0x1e7: frame_vm_group_bin_2178 (RW)
0x1e8: frame_vm_group_bin_18272 (RW)
0x1e9: frame_vm_group_bin_11184 (RW)
0x1e: frame_vm_group_bin_15396 (RW)
0x1ea: frame_vm_group_bin_3999 (RW)
0x1eb: frame_vm_group_bin_20096 (RW)
0x1ec: frame_vm_group_bin_12896 (RW)
0x1ed: frame_vm_group_bin_5804 (RW)
0x1ee: frame_vm_group_bin_21932 (RW)
0x1ef: frame_vm_group_bin_14757 (RW)
0x1f0: frame_vm_group_bin_7542 (RW)
0x1f1: frame_vm_group_bin_0387 (RW)
0x1f2: frame_vm_group_bin_16572 (RW)
0x1f3: frame_vm_group_bin_9361 (RW)
0x1f4: frame_vm_group_bin_17189 (RW)
0x1f5: frame_vm_group_bin_18305 (RW)
0x1f6: frame_vm_group_bin_11217 (RW)
0x1f7: frame_vm_group_bin_4032 (RW)
0x1f8: frame_vm_group_bin_20128 (RW)
0x1f9: frame_vm_group_bin_9980 (RW)
0x1f: frame_vm_group_bin_8205 (RW)
0x1fa: frame_vm_group_bin_5827 (RW)
0x1fb: frame_vm_group_bin_21966 (RW)
0x1fc: frame_vm_group_bin_14790 (RW)
0x1fd: frame_vm_group_bin_7575 (RW)
0x1fe: frame_vm_group_bin_0417 (RW)
0x1ff: frame_vm_group_bin_16605 (RW)
0x20: frame_vm_group_bin_12278 (RW)
0x21: frame_vm_group_bin_17241 (RW)
0x22: frame_vm_group_bin_10035 (RW)
0x23: frame_vm_group_bin_2878 (RW)
0x24: frame_vm_group_bin_18950 (RW)
0x25: frame_vm_group_bin_11807 (RW)
0x26: frame_vm_group_bin_4681 (RW)
0x27: frame_vm_group_bin_20803 (RW)
0x28: frame_vm_group_bin_13604 (RW)
0x29: frame_vm_group_bin_6414 (RW)
0x2: frame_vm_group_bin_6318 (RW)
0x2a: frame_vm_group_bin_22611 (RW)
0x2b: frame_vm_group_bin_15429 (RW)
0x2c: frame_vm_group_bin_8238 (RW)
0x2d: frame_vm_group_bin_17025 (RW)
0x2e: frame_vm_group_bin_17274 (RW)
0x2f: frame_vm_group_bin_10068 (RW)
0x30: frame_vm_group_bin_2911 (RW)
0x31: frame_vm_group_bin_18981 (RW)
0x32: frame_vm_group_bin_11839 (RW)
0x33: frame_vm_group_bin_4713 (RW)
0x34: frame_vm_group_bin_20835 (RW)
0x35: frame_vm_group_bin_13637 (RW)
0x36: frame_vm_group_bin_6447 (RW)
0x37: frame_vm_group_bin_22644 (RW)
0x38: frame_vm_group_bin_15462 (RW)
0x39: frame_vm_group_bin_8270 (RW)
0x3: frame_vm_group_bin_22512 (RW)
0x3a: frame_vm_group_bin_1087 (RW)
0x3b: frame_vm_group_bin_17308 (RW)
0x3c: frame_vm_group_bin_10102 (RW)
0x3d: frame_vm_group_bin_2945 (RW)
0x3e: frame_vm_group_bin_19015 (RW)
0x3f: frame_vm_group_bin_11869 (RW)
0x40: frame_vm_group_bin_4746 (RW)
0x41: frame_vm_group_bin_11640 (RW)
0x42: frame_vm_group_bin_13670 (RW)
0x43: frame_vm_group_bin_6481 (RW)
0x44: frame_vm_group_bin_22678 (RW)
0x45: frame_vm_group_bin_15496 (RW)
0x46: frame_vm_group_bin_8304 (RW)
0x47: frame_vm_group_bin_1115 (RW)
0x48: frame_vm_group_bin_17341 (RW)
0x49: frame_vm_group_bin_10135 (RW)
0x4: frame_vm_group_bin_15329 (RW)
0x4a: frame_vm_group_bin_2978 (RW)
0x4b: frame_vm_group_bin_19048 (RW)
0x4c: frame_vm_group_bin_11893 (RW)
0x4d: frame_vm_group_bin_4779 (RW)
0x4e: frame_vm_group_bin_20887 (RW)
0x4f: frame_vm_group_bin_13703 (RW)
0x50: frame_vm_group_bin_6514 (RW)
0x51: frame_vm_group_bin_22711 (RW)
0x52: frame_vm_group_bin_15528 (RW)
0x53: frame_vm_group_bin_8337 (RW)
0x54: frame_vm_group_bin_1148 (RW)
0x55: frame_vm_group_bin_17373 (RW)
0x56: frame_vm_group_bin_10170 (RW)
0x57: frame_vm_group_bin_3011 (RW)
0x58: frame_vm_group_bin_19081 (RW)
0x59: frame_vm_group_bin_11919 (RW)
0x5: frame_vm_group_bin_8138 (RW)
0x5a: frame_vm_group_bin_22387 (RW)
0x5b: frame_vm_group_bin_20917 (RW)
0x5c: frame_vm_group_bin_13736 (RW)
0x5d: frame_vm_group_bin_6548 (RW)
0x5e: frame_vm_group_bin_16672 (RW)
0x5f: frame_vm_group_bin_15561 (RW)
0x60: frame_vm_group_bin_8371 (RW)
0x61: frame_vm_group_bin_1182 (RW)
0x62: frame_vm_group_bin_17404 (RW)
0x63: frame_vm_group_bin_10204 (RW)
0x64: frame_vm_group_bin_3045 (RW)
0x65: frame_vm_group_bin_19114 (RW)
0x66: frame_vm_group_bin_11950 (RW)
0x67: frame_vm_group_bin_4845 (RW)
0x68: frame_vm_group_bin_2301 (RW)
0x69: frame_vm_group_bin_13770 (RW)
0x6: frame_vm_group_bin_0984 (RW)
0x6a: frame_vm_group_bin_6581 (RW)
0x6b: frame_vm_group_bin_22777 (RW)
0x6c: frame_vm_group_bin_15594 (RW)
0x6d: frame_vm_group_bin_8404 (RW)
0x6e: frame_vm_group_bin_1215 (RW)
0x6f: frame_vm_group_bin_15581 (RW)
0x70: frame_vm_group_bin_10237 (RW)
0x71: frame_vm_group_bin_3078 (RW)
0x72: frame_vm_group_bin_19146 (RW)
0x73: frame_vm_group_bin_11983 (RW)
0x74: frame_vm_group_bin_4878 (RW)
0x75: frame_vm_group_bin_20971 (RW)
0x76: frame_vm_group_bin_13803 (RW)
0x77: frame_vm_group_bin_6614 (RW)
0x78: frame_vm_group_bin_22810 (RW)
0x79: frame_vm_group_bin_15627 (RW)
0x7: frame_vm_group_bin_17177 (RW)
0x7a: frame_vm_group_bin_8438 (RW)
0x7b: frame_vm_group_bin_21680 (RW)
0x7c: frame_vm_group_bin_17454 (RW)
0x7d: frame_vm_group_bin_10271 (RW)
0x7e: frame_vm_group_bin_3112 (RW)
0x7f: frame_vm_group_bin_19180 (RW)
0x80: frame_vm_group_bin_12015 (RW)
0x81: frame_vm_group_bin_4912 (RW)
0x82: frame_vm_group_bin_21005 (RW)
0x83: frame_vm_group_bin_13835 (RW)
0x84: frame_vm_group_bin_6648 (RW)
0x85: frame_vm_group_bin_22844 (RW)
0x86: frame_vm_group_bin_15661 (RW)
0x87: frame_vm_group_bin_8471 (RW)
0x88: frame_vm_group_bin_1279 (RW)
0x89: frame_vm_group_bin_17472 (RW)
0x8: frame_vm_group_bin_9968 (RW)
0x8a: frame_vm_group_bin_10304 (RW)
0x8b: frame_vm_group_bin_3144 (RW)
0x8c: frame_vm_group_bin_19213 (RW)
0x8d: frame_vm_group_bin_12045 (RW)
0x8e: frame_vm_group_bin_4943 (RW)
0x8f: frame_vm_group_bin_21038 (RW)
0x90: frame_vm_group_bin_14883 (RW)
0x91: frame_vm_group_bin_6681 (RW)
0x92: frame_vm_group_bin_22877 (RW)
0x93: frame_vm_group_bin_15694 (RW)
0x94: frame_vm_group_bin_8504 (RW)
0x95: frame_vm_group_bin_1312 (RW)
0x96: frame_vm_group_bin_17495 (RW)
0x97: frame_vm_group_bin_10337 (RW)
0x98: frame_vm_group_bin_3177 (RW)
0x99: frame_vm_group_bin_19246 (RW)
0x9: frame_vm_group_bin_2810 (RW)
0x9a: frame_vm_group_bin_12074 (RW)
0x9b: frame_vm_group_bin_4975 (RW)
0x9c: frame_vm_group_bin_21073 (RW)
0x9d: frame_vm_group_bin_13895 (RW)
0x9e: frame_vm_group_bin_6714 (RW)
0x9f: frame_vm_group_bin_22911 (RW)
0xa0: frame_vm_group_bin_15728 (RW)
0xa1: frame_vm_group_bin_8537 (RW)
0xa2: frame_vm_group_bin_1345 (RW)
0xa3: frame_vm_group_bin_17521 (RW)
0xa4: frame_vm_group_bin_10371 (RW)
0xa5: frame_vm_group_bin_3211 (RW)
0xa6: frame_vm_group_bin_19280 (RW)
0xa7: frame_vm_group_bin_12107 (RW)
0xa8: frame_vm_group_bin_5008 (RW)
0xa9: frame_vm_group_bin_21106 (RW)
0xa: frame_vm_group_bin_18884 (RW)
0xaa: frame_vm_group_bin_13928 (RW)
0xab: frame_vm_group_bin_6747 (RW)
0xac: frame_vm_group_bin_22944 (RW)
0xad: frame_vm_group_bin_15761 (RW)
0xae: frame_vm_group_bin_8568 (RW)
0xaf: frame_vm_group_bin_1379 (RW)
0xb0: frame_vm_group_bin_17546 (RW)
0xb1: frame_vm_group_bin_14153 (RW)
0xb2: frame_vm_group_bin_3243 (RW)
0xb3: frame_vm_group_bin_19313 (RW)
0xb4: frame_vm_group_bin_12139 (RW)
0xb5: frame_vm_group_bin_5041 (RW)
0xb6: frame_vm_group_bin_21139 (RW)
0xb7: frame_vm_group_bin_13961 (RW)
0xb8: frame_vm_group_bin_6779 (RW)
0xb9: frame_vm_group_bin_22976 (RW)
0xb: frame_vm_group_bin_11752 (RW)
0xba: frame_vm_group_bin_15795 (RW)
0xbb: frame_vm_group_bin_8601 (RW)
0xbc: frame_vm_group_bin_1413 (RW)
0xbd: frame_vm_group_bin_17569 (RW)
0xbe: frame_vm_group_bin_10427 (RW)
0xbf: frame_vm_group_bin_3277 (RW)
0xc0: frame_vm_group_bin_19347 (RW)
0xc1: frame_vm_group_bin_12170 (RW)
0xc2: frame_vm_group_bin_5076 (RW)
0xc3: frame_vm_group_bin_21172 (RW)
0xc4: frame_vm_group_bin_13995 (RW)
0xc5: frame_vm_group_bin_6812 (RW)
0xc6: frame_vm_group_bin_23009 (RW)
0xc7: frame_vm_group_bin_15826 (RW)
0xc8: frame_vm_group_bin_8634 (RW)
0xc9: frame_vm_group_bin_1446 (RW)
0xc: frame_vm_group_bin_17668 (RW)
0xca: frame_vm_group_bin_17592 (RW)
0xcb: frame_vm_group_bin_10457 (RW)
0xcc: frame_vm_group_bin_3310 (RW)
0xcd: frame_vm_group_bin_19380 (RW)
0xce: frame_vm_group_bin_12202 (RW)
0xcf: frame_vm_group_bin_5109 (RW)
0xd0: frame_vm_group_bin_21205 (RW)
0xd1: frame_vm_group_bin_14028 (RW)
0xd2: frame_vm_group_bin_13426 (RW)
0xd3: frame_vm_group_bin_23042 (RW)
0xd4: frame_vm_group_bin_15859 (RW)
0xd5: frame_vm_group_bin_8667 (RW)
0xd6: frame_vm_group_bin_1479 (RW)
0xd7: frame_vm_group_bin_17619 (RW)
0xd8: frame_vm_group_bin_10490 (RW)
0xd9: frame_vm_group_bin_3343 (RW)
0xd: frame_vm_group_bin_20736 (RW)
0xda: frame_vm_group_bin_19414 (RW)
0xdb: frame_vm_group_bin_12232 (RW)
0xdc: frame_vm_group_bin_5143 (RW)
0xdd: frame_vm_group_bin_21239 (RW)
0xde: frame_vm_group_bin_14062 (RW)
0xdf: frame_vm_group_bin_6869 (RW)
0xe0: frame_vm_group_bin_23076 (RW)
0xe1: frame_vm_group_bin_15893 (RW)
0xe2: frame_vm_group_bin_8702 (RW)
0xe3: frame_vm_group_bin_1513 (RW)
0xe4: frame_vm_group_bin_17653 (RW)
0xe5: frame_vm_group_bin_10523 (RW)
0xe6: frame_vm_group_bin_3376 (RW)
0xe7: frame_vm_group_bin_19444 (RW)
0xe8: frame_vm_group_bin_12265 (RW)
0xe9: frame_vm_group_bin_5176 (RW)
0xe: frame_vm_group_bin_13537 (RW)
0xea: frame_vm_group_bin_21272 (RW)
0xeb: frame_vm_group_bin_14095 (RW)
0xec: frame_vm_group_bin_22812 (RW)
0xed: frame_vm_group_bin_23109 (RW)
0xee: frame_vm_group_bin_15926 (RW)
0xef: frame_vm_group_bin_8735 (RW)
0xf0: frame_vm_group_bin_1546 (RW)
0xf1: frame_vm_group_bin_17684 (RW)
0xf2: frame_vm_group_bin_10556 (RW)
0xf3: frame_vm_group_bin_3405 (RW)
0xf4: frame_vm_group_bin_19476 (RW)
0xf5: frame_vm_group_bin_12298 (RW)
0xf6: frame_vm_group_bin_5209 (RW)
0xf7: frame_vm_group_bin_21305 (RW)
0xf8: frame_vm_group_bin_14128 (RW)
0xf9: frame_vm_group_bin_6918 (RW)
0xf: frame_vm_group_bin_6351 (RW)
0xfa: frame_vm_group_bin_23142 (RW)
0xfb: frame_vm_group_bin_15960 (RW)
0xfc: frame_vm_group_bin_8769 (RW)
0xfd: frame_vm_group_bin_1580 (RW)
0xfe: frame_vm_group_bin_17712 (RW)
0xff: frame_vm_group_bin_10590 (RW)
}
pt_vm_group_bin_0035 {
0x0: frame_vm_group_bin_22912 (RW)
0x100: frame_vm_group_bin_5634 (RW)
0x101: frame_vm_group_bin_21734 (RW)
0x102: frame_vm_group_bin_14560 (RW)
0x103: frame_vm_group_bin_7345 (RW)
0x104: frame_vm_group_bin_0218 (RW)
0x105: frame_vm_group_bin_16374 (RW)
0x106: frame_vm_group_bin_9197 (RW)
0x107: frame_vm_group_bin_2011 (RW)
0x108: frame_vm_group_bin_18107 (RW)
0x109: frame_vm_group_bin_11019 (RW)
0x10: frame_vm_group_bin_1380 (RW)
0x10a: frame_vm_group_bin_3834 (RW)
0x10b: frame_vm_group_bin_19932 (RW)
0x10c: frame_vm_group_bin_12734 (RW)
0x10d: frame_vm_group_bin_5667 (RW)
0x10e: frame_vm_group_bin_21767 (RW)
0x10f: frame_vm_group_bin_14593 (RW)
0x110: frame_vm_group_bin_7378 (RW)
0x111: frame_vm_group_bin_0243 (RW)
0x112: frame_vm_group_bin_16407 (RW)
0x113: frame_vm_group_bin_13449 (RW)
0x114: frame_vm_group_bin_2044 (RW)
0x115: frame_vm_group_bin_18140 (RW)
0x116: frame_vm_group_bin_11052 (RW)
0x117: frame_vm_group_bin_3867 (RW)
0x118: frame_vm_group_bin_19965 (RW)
0x119: frame_vm_group_bin_12764 (RW)
0x11: frame_vm_group_bin_17547 (RW)
0x11a: frame_vm_group_bin_5701 (RW)
0x11b: frame_vm_group_bin_21801 (RW)
0x11c: frame_vm_group_bin_14626 (RW)
0x11d: frame_vm_group_bin_7412 (RW)
0x11e: frame_vm_group_bin_0266 (RW)
0x11f: frame_vm_group_bin_16441 (RW)
0x120: frame_vm_group_bin_18097 (RW)
0x121: frame_vm_group_bin_2078 (RW)
0x122: frame_vm_group_bin_18174 (RW)
0x123: frame_vm_group_bin_11086 (RW)
0x124: frame_vm_group_bin_3901 (RW)
0x125: frame_vm_group_bin_19997 (RW)
0x126: frame_vm_group_bin_12798 (RW)
0x127: frame_vm_group_bin_5734 (RW)
0x128: frame_vm_group_bin_21834 (RW)
0x129: frame_vm_group_bin_14659 (RW)
0x12: frame_vm_group_bin_9094 (RW)
0x12a: frame_vm_group_bin_7445 (RW)
0x12b: frame_vm_group_bin_0293 (RW)
0x12c: frame_vm_group_bin_16474 (RW)
0x12d: frame_vm_group_bin_22835 (RW)
0x12e: frame_vm_group_bin_2111 (RW)
0x12f: frame_vm_group_bin_18206 (RW)
0x130: frame_vm_group_bin_11119 (RW)
0x131: frame_vm_group_bin_3934 (RW)
0x132: frame_vm_group_bin_20030 (RW)
0x133: frame_vm_group_bin_12830 (RW)
0x134: frame_vm_group_bin_12723 (RW)
0x135: frame_vm_group_bin_21867 (RW)
0x136: frame_vm_group_bin_14692 (RW)
0x137: frame_vm_group_bin_7478 (RW)
0x138: frame_vm_group_bin_0325 (RW)
0x139: frame_vm_group_bin_16507 (RW)
0x13: frame_vm_group_bin_3244 (RW)
0x13a: frame_vm_group_bin_9299 (RW)
0x13b: frame_vm_group_bin_2146 (RW)
0x13c: frame_vm_group_bin_18240 (RW)
0x13d: frame_vm_group_bin_11152 (RW)
0x13e: frame_vm_group_bin_3967 (RW)
0x13f: frame_vm_group_bin_20064 (RW)
0x140: frame_vm_group_bin_12864 (RW)
0x141: frame_vm_group_bin_17466 (RW)
0x142: frame_vm_group_bin_21901 (RW)
0x143: frame_vm_group_bin_14726 (RW)
0x144: frame_vm_group_bin_7511 (RW)
0x145: frame_vm_group_bin_0357 (RW)
0x146: frame_vm_group_bin_16541 (RW)
0x147: frame_vm_group_bin_9329 (RW)
0x148: frame_vm_group_bin_2179 (RW)
0x149: frame_vm_group_bin_18273 (RW)
0x14: frame_vm_group_bin_19314 (RW)
0x14a: frame_vm_group_bin_11185 (RW)
0x14b: frame_vm_group_bin_4000 (RW)
0x14c: frame_vm_group_bin_20097 (RW)
0x14d: frame_vm_group_bin_12897 (RW)
0x14e: frame_vm_group_bin_5805 (RW)
0x14f: frame_vm_group_bin_21933 (RW)
0x150: frame_vm_group_bin_14758 (RW)
0x151: frame_vm_group_bin_7543 (RW)
0x152: frame_vm_group_bin_0388 (RW)
0x153: frame_vm_group_bin_16573 (RW)
0x154: frame_vm_group_bin_9362 (RW)
0x155: frame_vm_group_bin_12032 (RW)
0x156: frame_vm_group_bin_18306 (RW)
0x157: frame_vm_group_bin_11218 (RW)
0x158: frame_vm_group_bin_4033 (RW)
0x159: frame_vm_group_bin_20129 (RW)
0x15: frame_vm_group_bin_12140 (RW)
0x15a: frame_vm_group_bin_12930 (RW)
0x15b: frame_vm_group_bin_5828 (RW)
0x15c: frame_vm_group_bin_21967 (RW)
0x15d: frame_vm_group_bin_14791 (RW)
0x15e: frame_vm_group_bin_7576 (RW)
0x15f: frame_vm_group_bin_21022 (RW)
0x160: frame_vm_group_bin_16606 (RW)
0x161: frame_vm_group_bin_9397 (RW)
0x162: frame_vm_group_bin_2238 (RW)
0x163: frame_vm_group_bin_18340 (RW)
0x164: frame_vm_group_bin_11252 (RW)
0x165: frame_vm_group_bin_4067 (RW)
0x166: frame_vm_group_bin_20162 (RW)
0x167: frame_vm_group_bin_12963 (RW)
0x168: frame_vm_group_bin_5852 (RW)
0x169: frame_vm_group_bin_22000 (RW)
0x16: frame_vm_group_bin_5042 (RW)
0x16a: frame_vm_group_bin_14824 (RW)
0x16b: frame_vm_group_bin_7609 (RW)
0x16c: frame_vm_group_bin_0449 (RW)
0x16d: frame_vm_group_bin_16639 (RW)
0x16e: frame_vm_group_bin_9430 (RW)
0x16f: frame_vm_group_bin_2270 (RW)
0x170: frame_vm_group_bin_18373 (RW)
0x171: frame_vm_group_bin_11285 (RW)
0x172: frame_vm_group_bin_4100 (RW)
0x173: frame_vm_group_bin_20194 (RW)
0x174: frame_vm_group_bin_12996 (RW)
0x175: frame_vm_group_bin_5878 (RW)
0x176: frame_vm_group_bin_11407 (RW)
0x177: frame_vm_group_bin_14857 (RW)
0x178: frame_vm_group_bin_7642 (RW)
0x179: frame_vm_group_bin_0482 (RW)
0x17: frame_vm_group_bin_21140 (RW)
0x17a: frame_vm_group_bin_16673 (RW)
0x17b: frame_vm_group_bin_9464 (RW)
0x17c: frame_vm_group_bin_2304 (RW)
0x17d: frame_vm_group_bin_1291 (RW)
0x17e: frame_vm_group_bin_11319 (RW)
0x17f: frame_vm_group_bin_4133 (RW)
0x180: frame_vm_group_bin_20228 (RW)
0x181: frame_vm_group_bin_13032 (RW)
0x182: frame_vm_group_bin_5905 (RW)
0x183: frame_vm_group_bin_16056 (RW)
0x184: frame_vm_group_bin_14891 (RW)
0x185: frame_vm_group_bin_7676 (RW)
0x186: frame_vm_group_bin_0515 (RW)
0x187: frame_vm_group_bin_16705 (RW)
0x188: frame_vm_group_bin_9497 (RW)
0x189: frame_vm_group_bin_2337 (RW)
0x18: frame_vm_group_bin_13962 (RW)
0x18a: frame_vm_group_bin_18438 (RW)
0x18b: frame_vm_group_bin_11350 (RW)
0x18c: frame_vm_group_bin_4165 (RW)
0x18d: frame_vm_group_bin_20261 (RW)
0x18e: frame_vm_group_bin_13065 (RW)
0x18f: frame_vm_group_bin_5930 (RW)
0x190: frame_vm_group_bin_22075 (RW)
0x191: frame_vm_group_bin_14924 (RW)
0x192: frame_vm_group_bin_7709 (RW)
0x193: frame_vm_group_bin_0547 (RW)
0x194: frame_vm_group_bin_16739 (RW)
0x195: frame_vm_group_bin_9530 (RW)
0x196: frame_vm_group_bin_2370 (RW)
0x197: frame_vm_group_bin_18469 (RW)
0x198: frame_vm_group_bin_11382 (RW)
0x199: frame_vm_group_bin_4197 (RW)
0x19: frame_vm_group_bin_6780 (RW)
0x19a: frame_vm_group_bin_20294 (RW)
0x19b: frame_vm_group_bin_13099 (RW)
0x19c: frame_vm_group_bin_5952 (RW)
0x19d: frame_vm_group_bin_22107 (RW)
0x19e: frame_vm_group_bin_14958 (RW)
0x19f: frame_vm_group_bin_7742 (RW)
0x1: frame_vm_group_bin_15729 (RW)
0x1a0: frame_vm_group_bin_0579 (RW)
0x1a1: frame_vm_group_bin_16773 (RW)
0x1a2: frame_vm_group_bin_9564 (RW)
0x1a3: frame_vm_group_bin_2404 (RW)
0x1a4: frame_vm_group_bin_15321 (RW)
0x1a5: frame_vm_group_bin_11415 (RW)
0x1a6: frame_vm_group_bin_4231 (RW)
0x1a7: frame_vm_group_bin_20329 (RW)
0x1a8: frame_vm_group_bin_13132 (RW)
0x1a9: frame_vm_group_bin_5979 (RW)
0x1a: frame_vm_group_bin_22978 (RW)
0x1aa: frame_vm_group_bin_22140 (RW)
0x1ab: frame_vm_group_bin_14991 (RW)
0x1ac: frame_vm_group_bin_7775 (RW)
0x1ad: frame_vm_group_bin_0611 (RW)
0x1ae: frame_vm_group_bin_16806 (RW)
0x1af: frame_vm_group_bin_9597 (RW)
0x1b0: frame_vm_group_bin_2436 (RW)
0x1b1: frame_vm_group_bin_19967 (RW)
0x1b2: frame_vm_group_bin_11448 (RW)
0x1b3: frame_vm_group_bin_4264 (RW)
0x1b4: frame_vm_group_bin_20362 (RW)
0x1b5: frame_vm_group_bin_13165 (RW)
0x1b6: frame_vm_group_bin_6010 (RW)
0x1b7: frame_vm_group_bin_22173 (RW)
0x1b8: frame_vm_group_bin_15024 (RW)
0x1b9: frame_vm_group_bin_7808 (RW)
0x1b: frame_vm_group_bin_15796 (RW)
0x1ba: frame_vm_group_bin_0644 (RW)
0x1bb: frame_vm_group_bin_16840 (RW)
0x1bc: frame_vm_group_bin_9631 (RW)
0x1bd: frame_vm_group_bin_2469 (RW)
0x1be: frame_vm_group_bin_18550 (RW)
0x1bf: frame_vm_group_bin_11482 (RW)
0x1c0: frame_vm_group_bin_4298 (RW)
0x1c1: frame_vm_group_bin_20396 (RW)
0x1c2: frame_vm_group_bin_13199 (RW)
0x1c3: frame_vm_group_bin_6041 (RW)
0x1c4: frame_vm_group_bin_22207 (RW)
0x1c5: frame_vm_group_bin_14623 (RW)
0x1c6: frame_vm_group_bin_7841 (RW)
0x1c7: frame_vm_group_bin_0677 (RW)
0x1c8: frame_vm_group_bin_16872 (RW)
0x1c9: frame_vm_group_bin_9664 (RW)
0x1c: frame_vm_group_bin_8602 (RW)
0x1ca: frame_vm_group_bin_2502 (RW)
0x1cb: frame_vm_group_bin_18579 (RW)
0x1cc: frame_vm_group_bin_11515 (RW)
0x1cd: frame_vm_group_bin_4331 (RW)
0x1ce: frame_vm_group_bin_20429 (RW)
0x1cf: frame_vm_group_bin_13232 (RW)
0x1d0: frame_vm_group_bin_6064 (RW)
0x1d1: frame_vm_group_bin_22240 (RW)
0x1d2: frame_vm_group_bin_19247 (RW)
0x1d3: frame_vm_group_bin_7874 (RW)
0x1d4: frame_vm_group_bin_0710 (RW)
0x1d5: frame_vm_group_bin_16904 (RW)
0x1d6: frame_vm_group_bin_9696 (RW)
0x1d7: frame_vm_group_bin_2535 (RW)
0x1d8: frame_vm_group_bin_18612 (RW)
0x1d9: frame_vm_group_bin_11548 (RW)
0x1d: frame_vm_group_bin_1414 (RW)
0x1da: frame_vm_group_bin_4367 (RW)
0x1db: frame_vm_group_bin_20463 (RW)
0x1dc: frame_vm_group_bin_13266 (RW)
0x1dd: frame_vm_group_bin_6093 (RW)
0x1de: frame_vm_group_bin_22273 (RW)
0x1df: frame_vm_group_bin_15102 (RW)
0x1e0: frame_vm_group_bin_7908 (RW)
0x1e1: frame_vm_group_bin_0744 (RW)
0x1e2: frame_vm_group_bin_16938 (RW)
0x1e3: frame_vm_group_bin_9730 (RW)
0x1e4: frame_vm_group_bin_2569 (RW)
0x1e5: frame_vm_group_bin_18645 (RW)
0x1e6: frame_vm_group_bin_13891 (RW)
0x1e7: frame_vm_group_bin_4400 (RW)
0x1e8: frame_vm_group_bin_20496 (RW)
0x1e9: frame_vm_group_bin_13299 (RW)
0x1e: frame_vm_group_bin_17570 (RW)
0x1ea: frame_vm_group_bin_6124 (RW)
0x1eb: frame_vm_group_bin_22306 (RW)
0x1ec: frame_vm_group_bin_5352 (RW)
0x1ed: frame_vm_group_bin_7942 (RW)
0x1ee: frame_vm_group_bin_0777 (RW)
0x1ef: frame_vm_group_bin_16971 (RW)
0x1f0: frame_vm_group_bin_9763 (RW)
0x1f1: frame_vm_group_bin_2602 (RW)
0x1f2: frame_vm_group_bin_18678 (RW)
0x1f3: frame_vm_group_bin_18528 (RW)
0x1f4: frame_vm_group_bin_4433 (RW)
0x1f5: frame_vm_group_bin_20529 (RW)
0x1f6: frame_vm_group_bin_13331 (RW)
0x1f7: frame_vm_group_bin_6156 (RW)
0x1f8: frame_vm_group_bin_11453 (RW)
0x1f9: frame_vm_group_bin_15154 (RW)
0x1f: frame_vm_group_bin_10428 (RW)
0x1fa: frame_vm_group_bin_7976 (RW)
0x1fb: frame_vm_group_bin_0810 (RW)
0x1fc: frame_vm_group_bin_17005 (RW)
0x1fd: frame_vm_group_bin_9797 (RW)
0x1fe: frame_vm_group_bin_2636 (RW)
0x1ff: frame_vm_group_bin_18711 (RW)
0x20: frame_vm_group_bin_3278 (RW)
0x21: frame_vm_group_bin_19348 (RW)
0x22: frame_vm_group_bin_12171 (RW)
0x23: frame_vm_group_bin_5077 (RW)
0x24: frame_vm_group_bin_21173 (RW)
0x25: frame_vm_group_bin_13996 (RW)
0x26: frame_vm_group_bin_6813 (RW)
0x27: frame_vm_group_bin_23010 (RW)
0x28: frame_vm_group_bin_15827 (RW)
0x29: frame_vm_group_bin_8635 (RW)
0x2: frame_vm_group_bin_8538 (RW)
0x2a: frame_vm_group_bin_1447 (RW)
0x2b: frame_vm_group_bin_17593 (RW)
0x2c: frame_vm_group_bin_10458 (RW)
0x2d: frame_vm_group_bin_3311 (RW)
0x2e: frame_vm_group_bin_19381 (RW)
0x2f: frame_vm_group_bin_12203 (RW)
0x30: frame_vm_group_bin_5110 (RW)
0x31: frame_vm_group_bin_21206 (RW)
0x32: frame_vm_group_bin_14029 (RW)
0x33: frame_vm_group_bin_8366 (RW)
0x34: frame_vm_group_bin_23043 (RW)
0x35: frame_vm_group_bin_15860 (RW)
0x36: frame_vm_group_bin_8668 (RW)
0x37: frame_vm_group_bin_1480 (RW)
0x38: frame_vm_group_bin_17620 (RW)
0x39: frame_vm_group_bin_10491 (RW)
0x3: frame_vm_group_bin_1346 (RW)
0x3a: frame_vm_group_bin_3345 (RW)
0x3b: frame_vm_group_bin_20198 (RW)
0x3c: frame_vm_group_bin_12233 (RW)
0x3d: frame_vm_group_bin_5144 (RW)
0x3e: frame_vm_group_bin_21240 (RW)
0x3f: frame_vm_group_bin_14063 (RW)
0x40: frame_vm_group_bin_13001 (RW)
0x41: frame_vm_group_bin_23077 (RW)
0x42: frame_vm_group_bin_15894 (RW)
0x43: frame_vm_group_bin_8703 (RW)
0x44: frame_vm_group_bin_1514 (RW)
0x45: frame_vm_group_bin_17654 (RW)
0x46: frame_vm_group_bin_10524 (RW)
0x47: frame_vm_group_bin_3377 (RW)
0x48: frame_vm_group_bin_19445 (RW)
0x49: frame_vm_group_bin_12266 (RW)
0x4: frame_vm_group_bin_17522 (RW)
0x4a: frame_vm_group_bin_5177 (RW)
0x4b: frame_vm_group_bin_21273 (RW)
0x4c: frame_vm_group_bin_14096 (RW)
0x4d: frame_vm_group_bin_17689 (RW)
0x4e: frame_vm_group_bin_23110 (RW)
0x4f: frame_vm_group_bin_15927 (RW)
0x50: frame_vm_group_bin_8736 (RW)
0x51: frame_vm_group_bin_1547 (RW)
0x52: frame_vm_group_bin_17685 (RW)
0x53: frame_vm_group_bin_10557 (RW)
0x54: frame_vm_group_bin_7644 (RW)
0x55: frame_vm_group_bin_19477 (RW)
0x56: frame_vm_group_bin_12299 (RW)
0x57: frame_vm_group_bin_5210 (RW)
0x58: frame_vm_group_bin_1931 (RW)
0x59: frame_vm_group_bin_14129 (RW)
0x5: frame_vm_group_bin_10372 (RW)
0x5a: frame_vm_group_bin_6920 (RW)
0x5b: frame_vm_group_bin_23143 (RW)
0x5c: frame_vm_group_bin_15961 (RW)
0x5d: frame_vm_group_bin_8770 (RW)
0x5e: frame_vm_group_bin_1581 (RW)
0x5f: frame_vm_group_bin_17713 (RW)
0x60: frame_vm_group_bin_10591 (RW)
0x61: frame_vm_group_bin_12302 (RW)
0x62: frame_vm_group_bin_19511 (RW)
0x63: frame_vm_group_bin_12332 (RW)
0x64: frame_vm_group_bin_5244 (RW)
0x65: frame_vm_group_bin_21338 (RW)
0x66: frame_vm_group_bin_14163 (RW)
0x67: frame_vm_group_bin_6950 (RW)
0x68: frame_vm_group_bin_23176 (RW)
0x69: frame_vm_group_bin_15996 (RW)
0x6: frame_vm_group_bin_3212 (RW)
0x6a: frame_vm_group_bin_8803 (RW)
0x6b: frame_vm_group_bin_1614 (RW)
0x6c: frame_vm_group_bin_17739 (RW)
0x6d: frame_vm_group_bin_10624 (RW)
0x6e: frame_vm_group_bin_3451 (RW)
0x6f: frame_vm_group_bin_19544 (RW)
0x70: frame_vm_group_bin_12365 (RW)
0x71: frame_vm_group_bin_5277 (RW)
0x72: frame_vm_group_bin_21371 (RW)
0x73: frame_vm_group_bin_14195 (RW)
0x74: frame_vm_group_bin_6982 (RW)
0x75: frame_vm_group_bin_21798 (RW)
0x76: frame_vm_group_bin_16029 (RW)
0x77: frame_vm_group_bin_8836 (RW)
0x78: frame_vm_group_bin_1647 (RW)
0x79: frame_vm_group_bin_17767 (RW)
0x7: frame_vm_group_bin_19281 (RW)
0x7a: frame_vm_group_bin_23141 (RW)
0x7b: frame_vm_group_bin_3480 (RW)
0x7c: frame_vm_group_bin_19579 (RW)
0x7d: frame_vm_group_bin_12399 (RW)
0x7e: frame_vm_group_bin_17416 (RW)
0x7f: frame_vm_group_bin_21405 (RW)
0x80: frame_vm_group_bin_14229 (RW)
0x81: frame_vm_group_bin_7016 (RW)
0x82: frame_vm_group_bin_11657 (RW)
0x83: frame_vm_group_bin_16063 (RW)
0x84: frame_vm_group_bin_8869 (RW)
0x85: frame_vm_group_bin_1681 (RW)
0x86: frame_vm_group_bin_17798 (RW)
0x87: frame_vm_group_bin_10689 (RW)
0x88: frame_vm_group_bin_3506 (RW)
0x89: frame_vm_group_bin_19612 (RW)
0x8: frame_vm_group_bin_12108 (RW)
0x8a: frame_vm_group_bin_12432 (RW)
0x8b: frame_vm_group_bin_5342 (RW)
0x8c: frame_vm_group_bin_21437 (RW)
0x8d: frame_vm_group_bin_14261 (RW)
0x8e: frame_vm_group_bin_7048 (RW)
0x8f: frame_vm_group_bin_16319 (RW)
0x90: frame_vm_group_bin_16095 (RW)
0x91: frame_vm_group_bin_8901 (RW)
0x92: frame_vm_group_bin_1713 (RW)
0x93: frame_vm_group_bin_17828 (RW)
0x94: frame_vm_group_bin_10721 (RW)
0x95: frame_vm_group_bin_3535 (RW)
0x96: frame_vm_group_bin_19643 (RW)
0x97: frame_vm_group_bin_12463 (RW)
0x98: frame_vm_group_bin_5373 (RW)
0x99: frame_vm_group_bin_21469 (RW)
0x9: frame_vm_group_bin_5009 (RW)
0x9a: frame_vm_group_bin_14293 (RW)
0x9b: frame_vm_group_bin_7080 (RW)
0x9c: frame_vm_group_bin_0018 (RW)
0x9d: frame_vm_group_bin_16128 (RW)
0x9e: frame_vm_group_bin_8934 (RW)
0x9f: frame_vm_group_bin_1746 (RW)
0xa0: frame_vm_group_bin_17855 (RW)
0xa1: frame_vm_group_bin_10754 (RW)
0xa2: frame_vm_group_bin_3567 (RW)
0xa3: frame_vm_group_bin_19671 (RW)
0xa4: frame_vm_group_bin_12496 (RW)
0xa5: frame_vm_group_bin_5406 (RW)
0xa6: frame_vm_group_bin_21501 (RW)
0xa7: frame_vm_group_bin_14325 (RW)
0xa8: frame_vm_group_bin_7111 (RW)
0xa9: frame_vm_group_bin_0036 (RW)
0xa: frame_vm_group_bin_21107 (RW)
0xaa: frame_vm_group_bin_16159 (RW)
0xab: frame_vm_group_bin_8966 (RW)
0xac: frame_vm_group_bin_1778 (RW)
0xad: frame_vm_group_bin_17882 (RW)
0xae: frame_vm_group_bin_10786 (RW)
0xaf: frame_vm_group_bin_3601 (RW)
0xb0: frame_vm_group_bin_19701 (RW)
0xb1: frame_vm_group_bin_12529 (RW)
0xb2: frame_vm_group_bin_5439 (RW)
0xb3: frame_vm_group_bin_21534 (RW)
0xb4: frame_vm_group_bin_14358 (RW)
0xb5: frame_vm_group_bin_7143 (RW)
0xb6: frame_vm_group_bin_0061 (RW)
0xb7: frame_vm_group_bin_16192 (RW)
0xb8: frame_vm_group_bin_8999 (RW)
0xb9: frame_vm_group_bin_1811 (RW)
0xb: frame_vm_group_bin_13929 (RW)
0xba: frame_vm_group_bin_17914 (RW)
0xbb: frame_vm_group_bin_10820 (RW)
0xbc: frame_vm_group_bin_3635 (RW)
0xbd: frame_vm_group_bin_19735 (RW)
0xbe: frame_vm_group_bin_12563 (RW)
0xbf: frame_vm_group_bin_5471 (RW)
0xc0: frame_vm_group_bin_21568 (RW)
0xc1: frame_vm_group_bin_14392 (RW)
0xc2: frame_vm_group_bin_7179 (RW)
0xc3: frame_vm_group_bin_0088 (RW)
0xc4: frame_vm_group_bin_10244 (RW)
0xc5: frame_vm_group_bin_9033 (RW)
0xc6: frame_vm_group_bin_1845 (RW)
0xc7: frame_vm_group_bin_17946 (RW)
0xc8: frame_vm_group_bin_10853 (RW)
0xc9: frame_vm_group_bin_3668 (RW)
0xc: frame_vm_group_bin_6748 (RW)
0xca: frame_vm_group_bin_19768 (RW)
0xcb: frame_vm_group_bin_12596 (RW)
0xcc: frame_vm_group_bin_5504 (RW)
0xcd: frame_vm_group_bin_21601 (RW)
0xce: frame_vm_group_bin_14425 (RW)
0xcf: frame_vm_group_bin_7212 (RW)
0xd0: frame_vm_group_bin_0113 (RW)
0xd1: frame_vm_group_bin_14907 (RW)
0xd2: frame_vm_group_bin_9066 (RW)
0xd3: frame_vm_group_bin_1878 (RW)
0xd4: frame_vm_group_bin_17976 (RW)
0xd5: frame_vm_group_bin_10885 (RW)
0xd6: frame_vm_group_bin_3701 (RW)
0xd7: frame_vm_group_bin_19801 (RW)
0xd8: frame_vm_group_bin_12629 (RW)
0xd9: frame_vm_group_bin_5536 (RW)
0xd: frame_vm_group_bin_22945 (RW)
0xda: frame_vm_group_bin_21635 (RW)
0xdb: frame_vm_group_bin_14459 (RW)
0xdc: frame_vm_group_bin_7246 (RW)
0xdd: frame_vm_group_bin_0136 (RW)
0xde: frame_vm_group_bin_16277 (RW)
0xdf: frame_vm_group_bin_9100 (RW)
0xe0: frame_vm_group_bin_1912 (RW)
0xe1: frame_vm_group_bin_18010 (RW)
0xe2: frame_vm_group_bin_10920 (RW)
0xe3: frame_vm_group_bin_3735 (RW)
0xe4: frame_vm_group_bin_19835 (RW)
0xe5: frame_vm_group_bin_9509 (RW)
0xe6: frame_vm_group_bin_5570 (RW)
0xe7: frame_vm_group_bin_21668 (RW)
0xe8: frame_vm_group_bin_14492 (RW)
0xe9: frame_vm_group_bin_7279 (RW)
0xe: frame_vm_group_bin_15762 (RW)
0xea: frame_vm_group_bin_0157 (RW)
0xeb: frame_vm_group_bin_16308 (RW)
0xec: frame_vm_group_bin_9133 (RW)
0xed: frame_vm_group_bin_1945 (RW)
0xee: frame_vm_group_bin_18043 (RW)
0xef: frame_vm_group_bin_10953 (RW)
0xf0: frame_vm_group_bin_3768 (RW)
0xf1: frame_vm_group_bin_19868 (RW)
0xf2: frame_vm_group_bin_14176 (RW)
0xf3: frame_vm_group_bin_5602 (RW)
0xf4: frame_vm_group_bin_21700 (RW)
0xf5: frame_vm_group_bin_14526 (RW)
0xf6: frame_vm_group_bin_7311 (RW)
0xf7: frame_vm_group_bin_0186 (RW)
0xf8: frame_vm_group_bin_16340 (RW)
0xf9: frame_vm_group_bin_9164 (RW)
0xf: frame_vm_group_bin_8569 (RW)
0xfa: frame_vm_group_bin_1978 (RW)
0xfb: frame_vm_group_bin_18076 (RW)
0xfc: frame_vm_group_bin_10986 (RW)
0xfd: frame_vm_group_bin_3801 (RW)
0xfe: frame_vm_group_bin_19900 (RW)
0xff: frame_vm_group_bin_12710 (RW)
}
pt_vm_group_bin_0037 {
0x0: frame_vm_group_bin_13008 (RW)
0x100: frame_vm_group_bin_19017 (RW)
0x101: frame_vm_group_bin_11871 (RW)
0x102: frame_vm_group_bin_4748 (RW)
0x103: frame_vm_group_bin_1433 (RW)
0x104: frame_vm_group_bin_13672 (RW)
0x105: frame_vm_group_bin_6483 (RW)
0x106: frame_vm_group_bin_22680 (RW)
0x107: frame_vm_group_bin_15498 (RW)
0x108: frame_vm_group_bin_8306 (RW)
0x109: frame_vm_group_bin_1117 (RW)
0x10: frame_vm_group_bin_14900 (RW)
0x10a: frame_vm_group_bin_17343 (RW)
0x10b: frame_vm_group_bin_10137 (RW)
0x10c: frame_vm_group_bin_2980 (RW)
0x10d: frame_vm_group_bin_19050 (RW)
0x10e: frame_vm_group_bin_11895 (RW)
0x10f: frame_vm_group_bin_4781 (RW)
0x110: frame_vm_group_bin_20889 (RW)
0x111: frame_vm_group_bin_13705 (RW)
0x112: frame_vm_group_bin_6516 (RW)
0x113: frame_vm_group_bin_22713 (RW)
0x114: frame_vm_group_bin_15530 (RW)
0x115: frame_vm_group_bin_8339 (RW)
0x116: frame_vm_group_bin_1150 (RW)
0x117: frame_vm_group_bin_17375 (RW)
0x118: frame_vm_group_bin_10172 (RW)
0x119: frame_vm_group_bin_3013 (RW)
0x11: frame_vm_group_bin_7685 (RW)
0x11a: frame_vm_group_bin_19084 (RW)
0x11b: frame_vm_group_bin_11922 (RW)
0x11c: frame_vm_group_bin_4814 (RW)
0x11d: frame_vm_group_bin_10818 (RW)
0x11e: frame_vm_group_bin_13738 (RW)
0x11f: frame_vm_group_bin_6550 (RW)
0x120: frame_vm_group_bin_22746 (RW)
0x121: frame_vm_group_bin_15563 (RW)
0x122: frame_vm_group_bin_8373 (RW)
0x123: frame_vm_group_bin_1184 (RW)
0x124: frame_vm_group_bin_0738 (RW)
0x125: frame_vm_group_bin_10206 (RW)
0x126: frame_vm_group_bin_3047 (RW)
0x127: frame_vm_group_bin_19116 (RW)
0x128: frame_vm_group_bin_11952 (RW)
0x129: frame_vm_group_bin_4847 (RW)
0x12: frame_vm_group_bin_0524 (RW)
0x12a: frame_vm_group_bin_20945 (RW)
0x12b: frame_vm_group_bin_13772 (RW)
0x12c: frame_vm_group_bin_6583 (RW)
0x12d: frame_vm_group_bin_22779 (RW)
0x12e: frame_vm_group_bin_15596 (RW)
0x12f: frame_vm_group_bin_8406 (RW)
0x130: frame_vm_group_bin_1217 (RW)
0x131: frame_vm_group_bin_17428 (RW)
0x132: frame_vm_group_bin_10239 (RW)
0x133: frame_vm_group_bin_3080 (RW)
0x134: frame_vm_group_bin_19148 (RW)
0x135: frame_vm_group_bin_11985 (RW)
0x136: frame_vm_group_bin_4880 (RW)
0x137: frame_vm_group_bin_20973 (RW)
0x138: frame_vm_group_bin_13805 (RW)
0x139: frame_vm_group_bin_6616 (RW)
0x13: frame_vm_group_bin_16714 (RW)
0x13a: frame_vm_group_bin_22813 (RW)
0x13b: frame_vm_group_bin_15630 (RW)
0x13c: frame_vm_group_bin_8440 (RW)
0x13d: frame_vm_group_bin_1250 (RW)
0x13e: frame_vm_group_bin_17456 (RW)
0x13f: frame_vm_group_bin_10273 (RW)
0x140: frame_vm_group_bin_3113 (RW)
0x141: frame_vm_group_bin_19182 (RW)
0x142: frame_vm_group_bin_12017 (RW)
0x143: frame_vm_group_bin_4914 (RW)
0x144: frame_vm_group_bin_21007 (RW)
0x145: frame_vm_group_bin_0083 (RW)
0x146: frame_vm_group_bin_6650 (RW)
0x147: frame_vm_group_bin_22846 (RW)
0x148: frame_vm_group_bin_15663 (RW)
0x149: frame_vm_group_bin_8473 (RW)
0x14: frame_vm_group_bin_9506 (RW)
0x14a: frame_vm_group_bin_1281 (RW)
0x14b: frame_vm_group_bin_17474 (RW)
0x14c: frame_vm_group_bin_10306 (RW)
0x14d: frame_vm_group_bin_3146 (RW)
0x14e: frame_vm_group_bin_19215 (RW)
0x14f: frame_vm_group_bin_12047 (RW)
0x150: frame_vm_group_bin_4945 (RW)
0x151: frame_vm_group_bin_21040 (RW)
0x152: frame_vm_group_bin_13864 (RW)
0x153: frame_vm_group_bin_6683 (RW)
0x154: frame_vm_group_bin_22879 (RW)
0x155: frame_vm_group_bin_15696 (RW)
0x156: frame_vm_group_bin_8506 (RW)
0x157: frame_vm_group_bin_1313 (RW)
0x158: frame_vm_group_bin_17497 (RW)
0x159: frame_vm_group_bin_10339 (RW)
0x15: frame_vm_group_bin_2346 (RW)
0x15a: frame_vm_group_bin_3180 (RW)
0x15b: frame_vm_group_bin_19249 (RW)
0x15c: frame_vm_group_bin_12076 (RW)
0x15d: frame_vm_group_bin_4977 (RW)
0x15e: frame_vm_group_bin_21075 (RW)
0x15f: frame_vm_group_bin_13897 (RW)
0x160: frame_vm_group_bin_6716 (RW)
0x161: frame_vm_group_bin_22913 (RW)
0x162: frame_vm_group_bin_15730 (RW)
0x163: frame_vm_group_bin_8539 (RW)
0x164: frame_vm_group_bin_1347 (RW)
0x165: frame_vm_group_bin_17523 (RW)
0x166: frame_vm_group_bin_10373 (RW)
0x167: frame_vm_group_bin_3213 (RW)
0x168: frame_vm_group_bin_19282 (RW)
0x169: frame_vm_group_bin_12109 (RW)
0x16: frame_vm_group_bin_18447 (RW)
0x16a: frame_vm_group_bin_5010 (RW)
0x16b: frame_vm_group_bin_21108 (RW)
0x16c: frame_vm_group_bin_13930 (RW)
0x16d: frame_vm_group_bin_6749 (RW)
0x16e: frame_vm_group_bin_22946 (RW)
0x16f: frame_vm_group_bin_15763 (RW)
0x170: frame_vm_group_bin_8570 (RW)
0x171: frame_vm_group_bin_1381 (RW)
0x172: frame_vm_group_bin_17548 (RW)
0x173: frame_vm_group_bin_10400 (RW)
0x174: frame_vm_group_bin_3245 (RW)
0x175: frame_vm_group_bin_19315 (RW)
0x176: frame_vm_group_bin_12141 (RW)
0x177: frame_vm_group_bin_5043 (RW)
0x178: frame_vm_group_bin_20130 (RW)
0x179: frame_vm_group_bin_13963 (RW)
0x17: frame_vm_group_bin_11359 (RW)
0x17a: frame_vm_group_bin_6782 (RW)
0x17b: frame_vm_group_bin_22979 (RW)
0x17c: frame_vm_group_bin_15797 (RW)
0x17d: frame_vm_group_bin_8603 (RW)
0x17e: frame_vm_group_bin_1415 (RW)
0x17f: frame_vm_group_bin_17571 (RW)
0x180: frame_vm_group_bin_10429 (RW)
0x181: frame_vm_group_bin_3279 (RW)
0x182: frame_vm_group_bin_19349 (RW)
0x183: frame_vm_group_bin_12172 (RW)
0x184: frame_vm_group_bin_5078 (RW)
0x185: frame_vm_group_bin_21174 (RW)
0x186: frame_vm_group_bin_13997 (RW)
0x187: frame_vm_group_bin_6814 (RW)
0x188: frame_vm_group_bin_23011 (RW)
0x189: frame_vm_group_bin_15828 (RW)
0x18: frame_vm_group_bin_4174 (RW)
0x18a: frame_vm_group_bin_8636 (RW)
0x18b: frame_vm_group_bin_1448 (RW)
0x18c: frame_vm_group_bin_17594 (RW)
0x18d: frame_vm_group_bin_10459 (RW)
0x18e: frame_vm_group_bin_3312 (RW)
0x18f: frame_vm_group_bin_19382 (RW)
0x190: frame_vm_group_bin_12204 (RW)
0x191: frame_vm_group_bin_5111 (RW)
0x192: frame_vm_group_bin_21207 (RW)
0x193: frame_vm_group_bin_14030 (RW)
0x194: frame_vm_group_bin_6841 (RW)
0x195: frame_vm_group_bin_23044 (RW)
0x196: frame_vm_group_bin_15861 (RW)
0x197: frame_vm_group_bin_8669 (RW)
0x198: frame_vm_group_bin_1481 (RW)
0x199: frame_vm_group_bin_17621 (RW)
0x19: frame_vm_group_bin_20269 (RW)
0x19a: frame_vm_group_bin_10493 (RW)
0x19b: frame_vm_group_bin_3346 (RW)
0x19c: frame_vm_group_bin_19415 (RW)
0x19d: frame_vm_group_bin_12234 (RW)
0x19e: frame_vm_group_bin_5145 (RW)
0x19f: frame_vm_group_bin_21241 (RW)
0x1: frame_vm_group_bin_5885 (RW)
0x1a0: frame_vm_group_bin_14064 (RW)
0x1a1: frame_vm_group_bin_6870 (RW)
0x1a2: frame_vm_group_bin_23078 (RW)
0x1a3: frame_vm_group_bin_15895 (RW)
0x1a4: frame_vm_group_bin_8704 (RW)
0x1a5: frame_vm_group_bin_1515 (RW)
0x1a6: frame_vm_group_bin_17655 (RW)
0x1a7: frame_vm_group_bin_10525 (RW)
0x1a8: frame_vm_group_bin_3378 (RW)
0x1a9: frame_vm_group_bin_19446 (RW)
0x1a: frame_vm_group_bin_13075 (RW)
0x1aa: frame_vm_group_bin_12267 (RW)
0x1ab: frame_vm_group_bin_5178 (RW)
0x1ac: frame_vm_group_bin_21274 (RW)
0x1ad: frame_vm_group_bin_14097 (RW)
0x1ae: frame_vm_group_bin_6893 (RW)
0x1af: frame_vm_group_bin_23111 (RW)
0x1b0: frame_vm_group_bin_15928 (RW)
0x1b1: frame_vm_group_bin_8737 (RW)
0x1b2: frame_vm_group_bin_1548 (RW)
0x1b3: frame_vm_group_bin_17686 (RW)
0x1b4: frame_vm_group_bin_10558 (RW)
0x1b5: frame_vm_group_bin_2608 (RW)
0x1b6: frame_vm_group_bin_19478 (RW)
0x1b7: frame_vm_group_bin_12300 (RW)
0x1b8: frame_vm_group_bin_5211 (RW)
0x1b9: frame_vm_group_bin_21306 (RW)
0x1b: frame_vm_group_bin_5937 (RW)
0x1ba: frame_vm_group_bin_14131 (RW)
0x1bb: frame_vm_group_bin_6921 (RW)
0x1bc: frame_vm_group_bin_23144 (RW)
0x1bd: frame_vm_group_bin_15962 (RW)
0x1be: frame_vm_group_bin_8771 (RW)
0x1bf: frame_vm_group_bin_1582 (RW)
0x1c0: frame_vm_group_bin_17714 (RW)
0x1c1: frame_vm_group_bin_10592 (RW)
0x1c2: frame_vm_group_bin_3430 (RW)
0x1c3: frame_vm_group_bin_19512 (RW)
0x1c4: frame_vm_group_bin_12333 (RW)
0x1c5: frame_vm_group_bin_5245 (RW)
0x1c6: frame_vm_group_bin_21339 (RW)
0x1c7: frame_vm_group_bin_14164 (RW)
0x1c8: frame_vm_group_bin_6951 (RW)
0x1c9: frame_vm_group_bin_23177 (RW)
0x1c: frame_vm_group_bin_22085 (RW)
0x1ca: frame_vm_group_bin_15997 (RW)
0x1cb: frame_vm_group_bin_8804 (RW)
0x1cc: frame_vm_group_bin_1615 (RW)
0x1cd: frame_vm_group_bin_17740 (RW)
0x1ce: frame_vm_group_bin_10625 (RW)
0x1cf: frame_vm_group_bin_3452 (RW)
0x1d0: frame_vm_group_bin_19545 (RW)
0x1d1: frame_vm_group_bin_12366 (RW)
0x1d2: frame_vm_group_bin_5278 (RW)
0x1d3: frame_vm_group_bin_21372 (RW)
0x1d4: frame_vm_group_bin_14196 (RW)
0x1d5: frame_vm_group_bin_6983 (RW)
0x1d6: frame_vm_group_bin_23207 (RW)
0x1d7: frame_vm_group_bin_16030 (RW)
0x1d8: frame_vm_group_bin_8837 (RW)
0x1d9: frame_vm_group_bin_1648 (RW)
0x1d: frame_vm_group_bin_14934 (RW)
0x1da: frame_vm_group_bin_17769 (RW)
0x1db: frame_vm_group_bin_10657 (RW)
0x1dc: frame_vm_group_bin_3481 (RW)
0x1dd: frame_vm_group_bin_19580 (RW)
0x1de: frame_vm_group_bin_12400 (RW)
0x1df: frame_vm_group_bin_5311 (RW)
0x1e0: frame_vm_group_bin_21406 (RW)
0x1e1: frame_vm_group_bin_14230 (RW)
0x1e2: frame_vm_group_bin_7017 (RW)
0x1e3: frame_vm_group_bin_23229 (RW)
0x1e4: frame_vm_group_bin_16064 (RW)
0x1e5: frame_vm_group_bin_8870 (RW)
0x1e6: frame_vm_group_bin_1682 (RW)
0x1e7: frame_vm_group_bin_17799 (RW)
0x1e8: frame_vm_group_bin_10690 (RW)
0x1e9: frame_vm_group_bin_3507 (RW)
0x1e: frame_vm_group_bin_7718 (RW)
0x1ea: frame_vm_group_bin_19613 (RW)
0x1eb: frame_vm_group_bin_12433 (RW)
0x1ec: frame_vm_group_bin_5343 (RW)
0x1ed: frame_vm_group_bin_21438 (RW)
0x1ee: frame_vm_group_bin_14262 (RW)
0x1ef: frame_vm_group_bin_7049 (RW)
0x1f0: frame_vm_group_bin_23250 (RW)
0x1f1: frame_vm_group_bin_16096 (RW)
0x1f2: frame_vm_group_bin_8902 (RW)
0x1f3: frame_vm_group_bin_1714 (RW)
0x1f4: frame_vm_group_bin_17829 (RW)
0x1f5: frame_vm_group_bin_10722 (RW)
0x1f6: frame_vm_group_bin_3536 (RW)
0x1f7: frame_vm_group_bin_19644 (RW)
0x1f8: frame_vm_group_bin_12464 (RW)
0x1f9: frame_vm_group_bin_5374 (RW)
0x1f: frame_vm_group_bin_0556 (RW)
0x1fa: frame_vm_group_bin_21471 (RW)
0x1fb: frame_vm_group_bin_14294 (RW)
0x1fc: frame_vm_group_bin_7081 (RW)
0x1fd: frame_vm_group_bin_0019 (RW)
0x1fe: frame_vm_group_bin_16129 (RW)
0x1ff: frame_vm_group_bin_8935 (RW)
0x20: frame_vm_group_bin_16749 (RW)
0x21: frame_vm_group_bin_9540 (RW)
0x22: frame_vm_group_bin_2380 (RW)
0x23: frame_vm_group_bin_19646 (RW)
0x24: frame_vm_group_bin_11392 (RW)
0x25: frame_vm_group_bin_4207 (RW)
0x26: frame_vm_group_bin_20303 (RW)
0x27: frame_vm_group_bin_13108 (RW)
0x28: frame_vm_group_bin_5959 (RW)
0x29: frame_vm_group_bin_22116 (RW)
0x2: frame_vm_group_bin_20365 (RW)
0x2a: frame_vm_group_bin_14967 (RW)
0x2b: frame_vm_group_bin_7751 (RW)
0x2c: frame_vm_group_bin_0587 (RW)
0x2d: frame_vm_group_bin_16782 (RW)
0x2e: frame_vm_group_bin_9573 (RW)
0x2f: frame_vm_group_bin_2413 (RW)
0x30: frame_vm_group_bin_18503 (RW)
0x31: frame_vm_group_bin_11424 (RW)
0x32: frame_vm_group_bin_4240 (RW)
0x33: frame_vm_group_bin_20338 (RW)
0x34: frame_vm_group_bin_13141 (RW)
0x35: frame_vm_group_bin_5988 (RW)
0x36: frame_vm_group_bin_22149 (RW)
0x37: frame_vm_group_bin_15000 (RW)
0x38: frame_vm_group_bin_7784 (RW)
0x39: frame_vm_group_bin_0620 (RW)
0x3: frame_vm_group_bin_14867 (RW)
0x3a: frame_vm_group_bin_16816 (RW)
0x3b: frame_vm_group_bin_9607 (RW)
0x3c: frame_vm_group_bin_2446 (RW)
0x3d: frame_vm_group_bin_18532 (RW)
0x3e: frame_vm_group_bin_11458 (RW)
0x3f: frame_vm_group_bin_4274 (RW)
0x40: frame_vm_group_bin_20372 (RW)
0x41: frame_vm_group_bin_13175 (RW)
0x42: frame_vm_group_bin_6019 (RW)
0x43: frame_vm_group_bin_22183 (RW)
0x44: frame_vm_group_bin_18920 (RW)
0x45: frame_vm_group_bin_7818 (RW)
0x46: frame_vm_group_bin_0653 (RW)
0x47: frame_vm_group_bin_16849 (RW)
0x48: frame_vm_group_bin_9640 (RW)
0x49: frame_vm_group_bin_2478 (RW)
0x4: frame_vm_group_bin_7652 (RW)
0x4a: frame_vm_group_bin_18557 (RW)
0x4b: frame_vm_group_bin_11491 (RW)
0x4c: frame_vm_group_bin_4307 (RW)
0x4d: frame_vm_group_bin_20405 (RW)
0x4e: frame_vm_group_bin_13208 (RW)
0x4f: frame_vm_group_bin_6047 (RW)
0x50: frame_vm_group_bin_22216 (RW)
0x51: frame_vm_group_bin_15057 (RW)
0x52: frame_vm_group_bin_7850 (RW)
0x53: frame_vm_group_bin_0686 (RW)
0x54: frame_vm_group_bin_16881 (RW)
0x55: frame_vm_group_bin_9673 (RW)
0x56: frame_vm_group_bin_2511 (RW)
0x57: frame_vm_group_bin_18588 (RW)
0x58: frame_vm_group_bin_11524 (RW)
0x59: frame_vm_group_bin_4342 (RW)
0x5: frame_vm_group_bin_0491 (RW)
0x5a: frame_vm_group_bin_20439 (RW)
0x5b: frame_vm_group_bin_13242 (RW)
0x5c: frame_vm_group_bin_6072 (RW)
0x5d: frame_vm_group_bin_22250 (RW)
0x5e: frame_vm_group_bin_15084 (RW)
0x5f: frame_vm_group_bin_7884 (RW)
0x60: frame_vm_group_bin_0720 (RW)
0x61: frame_vm_group_bin_16914 (RW)
0x62: frame_vm_group_bin_9706 (RW)
0x63: frame_vm_group_bin_2545 (RW)
0x64: frame_vm_group_bin_18622 (RW)
0x65: frame_vm_group_bin_3584 (RW)
0x66: frame_vm_group_bin_4376 (RW)
0x67: frame_vm_group_bin_20472 (RW)
0x68: frame_vm_group_bin_13275 (RW)
0x69: frame_vm_group_bin_6102 (RW)
0x6: frame_vm_group_bin_16682 (RW)
0x6a: frame_vm_group_bin_22282 (RW)
0x6b: frame_vm_group_bin_15108 (RW)
0x6c: frame_vm_group_bin_7917 (RW)
0x6d: frame_vm_group_bin_0753 (RW)
0x6e: frame_vm_group_bin_16947 (RW)
0x6f: frame_vm_group_bin_9739 (RW)
0x70: frame_vm_group_bin_2578 (RW)
0x71: frame_vm_group_bin_18654 (RW)
0x72: frame_vm_group_bin_22954 (RW)
0x73: frame_vm_group_bin_4409 (RW)
0x74: frame_vm_group_bin_20505 (RW)
0x75: frame_vm_group_bin_13308 (RW)
0x76: frame_vm_group_bin_6133 (RW)
0x77: frame_vm_group_bin_22315 (RW)
0x78: frame_vm_group_bin_15134 (RW)
0x79: frame_vm_group_bin_7951 (RW)
0x7: frame_vm_group_bin_9473 (RW)
0x7a: frame_vm_group_bin_0787 (RW)
0x7b: frame_vm_group_bin_16981 (RW)
0x7c: frame_vm_group_bin_9773 (RW)
0x7d: frame_vm_group_bin_2612 (RW)
0x7e: frame_vm_group_bin_18688 (RW)
0x7f: frame_vm_group_bin_11611 (RW)
0x80: frame_vm_group_bin_4443 (RW)
0x81: frame_vm_group_bin_20539 (RW)
0x82: frame_vm_group_bin_13341 (RW)
0x83: frame_vm_group_bin_6166 (RW)
0x84: frame_vm_group_bin_22348 (RW)
0x85: frame_vm_group_bin_15164 (RW)
0x86: frame_vm_group_bin_7985 (RW)
0x87: frame_vm_group_bin_0819 (RW)
0x88: frame_vm_group_bin_17014 (RW)
0x89: frame_vm_group_bin_9806 (RW)
0x8: frame_vm_group_bin_2313 (RW)
0x8a: frame_vm_group_bin_2645 (RW)
0x8b: frame_vm_group_bin_18720 (RW)
0x8c: frame_vm_group_bin_11633 (RW)
0x8d: frame_vm_group_bin_4476 (RW)
0x8e: frame_vm_group_bin_20572 (RW)
0x8f: frame_vm_group_bin_13373 (RW)
0x90: frame_vm_group_bin_6197 (RW)
0x91: frame_vm_group_bin_22381 (RW)
0x92: frame_vm_group_bin_15197 (RW)
0x93: frame_vm_group_bin_8014 (RW)
0x94: frame_vm_group_bin_0852 (RW)
0x95: frame_vm_group_bin_17047 (RW)
0x96: frame_vm_group_bin_9839 (RW)
0x97: frame_vm_group_bin_2678 (RW)
0x98: frame_vm_group_bin_18751 (RW)
0x99: frame_vm_group_bin_11656 (RW)
0x9: frame_vm_group_bin_18414 (RW)
0x9a: frame_vm_group_bin_4510 (RW)
0x9b: frame_vm_group_bin_20606 (RW)
0x9c: frame_vm_group_bin_13406 (RW)
0x9d: frame_vm_group_bin_6225 (RW)
0x9e: frame_vm_group_bin_6402 (RW)
0x9f: frame_vm_group_bin_15232 (RW)
0xa0: frame_vm_group_bin_8044 (RW)
0xa1: frame_vm_group_bin_0886 (RW)
0xa2: frame_vm_group_bin_17081 (RW)
0xa3: frame_vm_group_bin_9873 (RW)
0xa4: frame_vm_group_bin_2712 (RW)
0xa5: frame_vm_group_bin_18785 (RW)
0xa6: frame_vm_group_bin_11680 (RW)
0xa7: frame_vm_group_bin_4543 (RW)
0xa8: frame_vm_group_bin_20639 (RW)
0xa9: frame_vm_group_bin_13439 (RW)
0xa: frame_vm_group_bin_11328 (RW)
0xaa: frame_vm_group_bin_6255 (RW)
0xab: frame_vm_group_bin_22447 (RW)
0xac: frame_vm_group_bin_15265 (RW)
0xad: frame_vm_group_bin_8075 (RW)
0xae: frame_vm_group_bin_0919 (RW)
0xaf: frame_vm_group_bin_17114 (RW)
0xb0: frame_vm_group_bin_9905 (RW)
0xb1: frame_vm_group_bin_2745 (RW)
0xb2: frame_vm_group_bin_18818 (RW)
0xb3: frame_vm_group_bin_11707 (RW)
0xb4: frame_vm_group_bin_21515 (RW)
0xb5: frame_vm_group_bin_20671 (RW)
0xb6: frame_vm_group_bin_13472 (RW)
0xb7: frame_vm_group_bin_6287 (RW)
0xb8: frame_vm_group_bin_22480 (RW)
0xb9: frame_vm_group_bin_15297 (RW)
0xb: frame_vm_group_bin_4142 (RW)
0xba: frame_vm_group_bin_8108 (RW)
0xbb: frame_vm_group_bin_0953 (RW)
0xbc: frame_vm_group_bin_10052 (RW)
0xbd: frame_vm_group_bin_9937 (RW)
0xbe: frame_vm_group_bin_2779 (RW)
0xbf: frame_vm_group_bin_18853 (RW)
0xc0: frame_vm_group_bin_11733 (RW)
0xc1: frame_vm_group_bin_4596 (RW)
0xc2: frame_vm_group_bin_20705 (RW)
0xc3: frame_vm_group_bin_13506 (RW)
0xc4: frame_vm_group_bin_6320 (RW)
0xc5: frame_vm_group_bin_22514 (RW)
0xc6: frame_vm_group_bin_15331 (RW)
0xc7: frame_vm_group_bin_8140 (RW)
0xc8: frame_vm_group_bin_0986 (RW)
0xc9: frame_vm_group_bin_17179 (RW)
0xc: frame_vm_group_bin_20237 (RW)
0xca: frame_vm_group_bin_9970 (RW)
0xcb: frame_vm_group_bin_2812 (RW)
0xcc: frame_vm_group_bin_18886 (RW)
0xcd: frame_vm_group_bin_11754 (RW)
0xce: frame_vm_group_bin_4620 (RW)
0xcf: frame_vm_group_bin_20738 (RW)
0xd0: frame_vm_group_bin_13539 (RW)
0xd1: frame_vm_group_bin_6353 (RW)
0xd2: frame_vm_group_bin_22546 (RW)
0xd3: frame_vm_group_bin_15364 (RW)
0xd4: frame_vm_group_bin_8173 (RW)
0xd5: frame_vm_group_bin_20815 (RW)
0xd6: frame_vm_group_bin_17210 (RW)
0xd7: frame_vm_group_bin_10003 (RW)
0xd8: frame_vm_group_bin_2845 (RW)
0xd9: frame_vm_group_bin_18919 (RW)
0xd: frame_vm_group_bin_13041 (RW)
0xda: frame_vm_group_bin_11780 (RW)
0xdb: frame_vm_group_bin_4651 (RW)
0xdc: frame_vm_group_bin_20772 (RW)
0xdd: frame_vm_group_bin_13573 (RW)
0xde: frame_vm_group_bin_6384 (RW)
0xdf: frame_vm_group_bin_22580 (RW)
0xe0: frame_vm_group_bin_15398 (RW)
0xe1: frame_vm_group_bin_8207 (RW)
0xe2: frame_vm_group_bin_1041 (RW)
0xe3: frame_vm_group_bin_17243 (RW)
0xe4: frame_vm_group_bin_10037 (RW)
0xe5: frame_vm_group_bin_2880 (RW)
0xe6: frame_vm_group_bin_18952 (RW)
0xe7: frame_vm_group_bin_11809 (RW)
0xe8: frame_vm_group_bin_4683 (RW)
0xe9: frame_vm_group_bin_20805 (RW)
0xe: frame_vm_group_bin_5911 (RW)
0xea: frame_vm_group_bin_13606 (RW)
0xeb: frame_vm_group_bin_6416 (RW)
0xec: frame_vm_group_bin_22613 (RW)
0xed: frame_vm_group_bin_15431 (RW)
0xee: frame_vm_group_bin_8240 (RW)
0xef: frame_vm_group_bin_1061 (RW)
0xf0: frame_vm_group_bin_17276 (RW)
0xf1: frame_vm_group_bin_10070 (RW)
0xf2: frame_vm_group_bin_2913 (RW)
0xf3: frame_vm_group_bin_18983 (RW)
0xf4: frame_vm_group_bin_11841 (RW)
0xf5: frame_vm_group_bin_4715 (RW)
0xf6: frame_vm_group_bin_20837 (RW)
0xf7: frame_vm_group_bin_13638 (RW)
0xf8: frame_vm_group_bin_6449 (RW)
0xf9: frame_vm_group_bin_22646 (RW)
0xf: frame_vm_group_bin_22056 (RW)
0xfa: frame_vm_group_bin_15465 (RW)
0xfb: frame_vm_group_bin_8273 (RW)
0xfc: frame_vm_group_bin_1089 (RW)
0xfd: frame_vm_group_bin_17310 (RW)
0xfe: frame_vm_group_bin_10104 (RW)
0xff: frame_vm_group_bin_2947 (RW)
}
pt_vm_group_bin_0039 {
0x0: frame_vm_group_bin_15233 (RW)
0x100: frame_vm_group_bin_21242 (RW)
0x101: frame_vm_group_bin_14065 (RW)
0x102: frame_vm_group_bin_6871 (RW)
0x103: frame_vm_group_bin_23079 (RW)
0x104: frame_vm_group_bin_15896 (RW)
0x105: frame_vm_group_bin_8705 (RW)
0x106: frame_vm_group_bin_1516 (RW)
0x107: frame_vm_group_bin_17656 (RW)
0x108: frame_vm_group_bin_10526 (RW)
0x109: frame_vm_group_bin_16195 (RW)
0x10: frame_vm_group_bin_17115 (RW)
0x10a: frame_vm_group_bin_19447 (RW)
0x10b: frame_vm_group_bin_12268 (RW)
0x10c: frame_vm_group_bin_5179 (RW)
0x10d: frame_vm_group_bin_21275 (RW)
0x10e: frame_vm_group_bin_14098 (RW)
0x10f: frame_vm_group_bin_6894 (RW)
0x110: frame_vm_group_bin_23112 (RW)
0x111: frame_vm_group_bin_15929 (RW)
0x112: frame_vm_group_bin_8738 (RW)
0x113: frame_vm_group_bin_1549 (RW)
0x114: frame_vm_group_bin_17687 (RW)
0x115: frame_vm_group_bin_10559 (RW)
0x116: frame_vm_group_bin_20839 (RW)
0x117: frame_vm_group_bin_19479 (RW)
0x118: frame_vm_group_bin_12301 (RW)
0x119: frame_vm_group_bin_5212 (RW)
0x11: frame_vm_group_bin_9906 (RW)
0x11a: frame_vm_group_bin_21308 (RW)
0x11b: frame_vm_group_bin_14132 (RW)
0x11c: frame_vm_group_bin_6922 (RW)
0x11d: frame_vm_group_bin_23145 (RW)
0x11e: frame_vm_group_bin_15963 (RW)
0x11f: frame_vm_group_bin_8772 (RW)
0x120: frame_vm_group_bin_1583 (RW)
0x121: frame_vm_group_bin_17715 (RW)
0x122: frame_vm_group_bin_10593 (RW)
0x123: frame_vm_group_bin_3431 (RW)
0x124: frame_vm_group_bin_19513 (RW)
0x125: frame_vm_group_bin_12334 (RW)
0x126: frame_vm_group_bin_5246 (RW)
0x127: frame_vm_group_bin_21340 (RW)
0x128: frame_vm_group_bin_14165 (RW)
0x129: frame_vm_group_bin_6952 (RW)
0x12: frame_vm_group_bin_2746 (RW)
0x12a: frame_vm_group_bin_23178 (RW)
0x12b: frame_vm_group_bin_15998 (RW)
0x12c: frame_vm_group_bin_8805 (RW)
0x12d: frame_vm_group_bin_1616 (RW)
0x12e: frame_vm_group_bin_17741 (RW)
0x12f: frame_vm_group_bin_10626 (RW)
0x130: frame_vm_group_bin_3453 (RW)
0x131: frame_vm_group_bin_19546 (RW)
0x132: frame_vm_group_bin_12367 (RW)
0x133: frame_vm_group_bin_5279 (RW)
0x134: frame_vm_group_bin_21373 (RW)
0x135: frame_vm_group_bin_14197 (RW)
0x136: frame_vm_group_bin_6984 (RW)
0x137: frame_vm_group_bin_20107 (RW)
0x138: frame_vm_group_bin_16031 (RW)
0x139: frame_vm_group_bin_8838 (RW)
0x13: frame_vm_group_bin_18819 (RW)
0x13a: frame_vm_group_bin_1650 (RW)
0x13b: frame_vm_group_bin_17770 (RW)
0x13c: frame_vm_group_bin_10658 (RW)
0x13d: frame_vm_group_bin_3482 (RW)
0x13e: frame_vm_group_bin_19581 (RW)
0x13f: frame_vm_group_bin_12401 (RW)
0x140: frame_vm_group_bin_5312 (RW)
0x141: frame_vm_group_bin_21407 (RW)
0x142: frame_vm_group_bin_14231 (RW)
0x143: frame_vm_group_bin_7018 (RW)
0x144: frame_vm_group_bin_23230 (RW)
0x145: frame_vm_group_bin_16065 (RW)
0x146: frame_vm_group_bin_8871 (RW)
0x147: frame_vm_group_bin_1683 (RW)
0x148: frame_vm_group_bin_17800 (RW)
0x149: frame_vm_group_bin_10691 (RW)
0x14: frame_vm_group_bin_11708 (RW)
0x14a: frame_vm_group_bin_3508 (RW)
0x14b: frame_vm_group_bin_19614 (RW)
0x14c: frame_vm_group_bin_13286 (RW)
0x14d: frame_vm_group_bin_5344 (RW)
0x14e: frame_vm_group_bin_21439 (RW)
0x14f: frame_vm_group_bin_14263 (RW)
0x150: frame_vm_group_bin_7050 (RW)
0x151: frame_vm_group_bin_23251 (RW)
0x152: frame_vm_group_bin_16097 (RW)
0x153: frame_vm_group_bin_8903 (RW)
0x154: frame_vm_group_bin_1715 (RW)
0x155: frame_vm_group_bin_17830 (RW)
0x156: frame_vm_group_bin_10723 (RW)
0x157: frame_vm_group_bin_3537 (RW)
0x158: frame_vm_group_bin_19645 (RW)
0x159: frame_vm_group_bin_12465 (RW)
0x15: frame_vm_group_bin_16460 (RW)
0x15a: frame_vm_group_bin_5376 (RW)
0x15b: frame_vm_group_bin_21472 (RW)
0x15c: frame_vm_group_bin_14295 (RW)
0x15d: frame_vm_group_bin_7082 (RW)
0x15e: frame_vm_group_bin_0020 (RW)
0x15f: frame_vm_group_bin_9365 (RW)
0x160: frame_vm_group_bin_8936 (RW)
0x161: frame_vm_group_bin_1748 (RW)
0x162: frame_vm_group_bin_17857 (RW)
0x163: frame_vm_group_bin_10756 (RW)
0x164: frame_vm_group_bin_3569 (RW)
0x165: frame_vm_group_bin_19673 (RW)
0x166: frame_vm_group_bin_12498 (RW)
0x167: frame_vm_group_bin_5408 (RW)
0x168: frame_vm_group_bin_21503 (RW)
0x169: frame_vm_group_bin_14327 (RW)
0x16: frame_vm_group_bin_20672 (RW)
0x16a: frame_vm_group_bin_7113 (RW)
0x16b: frame_vm_group_bin_0038 (RW)
0x16c: frame_vm_group_bin_16161 (RW)
0x16d: frame_vm_group_bin_8968 (RW)
0x16e: frame_vm_group_bin_1780 (RW)
0x16f: frame_vm_group_bin_17884 (RW)
0x170: frame_vm_group_bin_10788 (RW)
0x171: frame_vm_group_bin_3603 (RW)
0x172: frame_vm_group_bin_19703 (RW)
0x173: frame_vm_group_bin_12531 (RW)
0x174: frame_vm_group_bin_5441 (RW)
0x175: frame_vm_group_bin_21536 (RW)
0x176: frame_vm_group_bin_14360 (RW)
0x177: frame_vm_group_bin_7145 (RW)
0x178: frame_vm_group_bin_0063 (RW)
0x179: frame_vm_group_bin_16194 (RW)
0x17: frame_vm_group_bin_13473 (RW)
0x17a: frame_vm_group_bin_9002 (RW)
0x17b: frame_vm_group_bin_1814 (RW)
0x17c: frame_vm_group_bin_17916 (RW)
0x17d: frame_vm_group_bin_10822 (RW)
0x17e: frame_vm_group_bin_3637 (RW)
0x17f: frame_vm_group_bin_19737 (RW)
0x180: frame_vm_group_bin_12565 (RW)
0x181: frame_vm_group_bin_5473 (RW)
0x182: frame_vm_group_bin_21570 (RW)
0x183: frame_vm_group_bin_14394 (RW)
0x184: frame_vm_group_bin_7181 (RW)
0x185: frame_vm_group_bin_0090 (RW)
0x186: frame_vm_group_bin_16222 (RW)
0x187: frame_vm_group_bin_9035 (RW)
0x188: frame_vm_group_bin_1847 (RW)
0x189: frame_vm_group_bin_17948 (RW)
0x18: frame_vm_group_bin_6288 (RW)
0x18a: frame_vm_group_bin_10855 (RW)
0x18b: frame_vm_group_bin_3670 (RW)
0x18c: frame_vm_group_bin_19770 (RW)
0x18d: frame_vm_group_bin_12598 (RW)
0x18e: frame_vm_group_bin_5506 (RW)
0x18f: frame_vm_group_bin_21603 (RW)
0x190: frame_vm_group_bin_14427 (RW)
0x191: frame_vm_group_bin_7214 (RW)
0x192: frame_vm_group_bin_0115 (RW)
0x193: frame_vm_group_bin_16248 (RW)
0x194: frame_vm_group_bin_9068 (RW)
0x195: frame_vm_group_bin_1880 (RW)
0x196: frame_vm_group_bin_17978 (RW)
0x197: frame_vm_group_bin_10887 (RW)
0x198: frame_vm_group_bin_3703 (RW)
0x199: frame_vm_group_bin_19803 (RW)
0x19: frame_vm_group_bin_22481 (RW)
0x19a: frame_vm_group_bin_12632 (RW)
0x19b: frame_vm_group_bin_5539 (RW)
0x19c: frame_vm_group_bin_21637 (RW)
0x19d: frame_vm_group_bin_14461 (RW)
0x19e: frame_vm_group_bin_7248 (RW)
0x19f: frame_vm_group_bin_0138 (RW)
0x1: frame_vm_group_bin_8045 (RW)
0x1a0: frame_vm_group_bin_16279 (RW)
0x1a1: frame_vm_group_bin_9102 (RW)
0x1a2: frame_vm_group_bin_1914 (RW)
0x1a3: frame_vm_group_bin_18012 (RW)
0x1a4: frame_vm_group_bin_10922 (RW)
0x1a5: frame_vm_group_bin_3737 (RW)
0x1a6: frame_vm_group_bin_19837 (RW)
0x1a7: frame_vm_group_bin_12661 (RW)
0x1a8: frame_vm_group_bin_5572 (RW)
0x1a9: frame_vm_group_bin_21670 (RW)
0x1a: frame_vm_group_bin_15299 (RW)
0x1aa: frame_vm_group_bin_14494 (RW)
0x1ab: frame_vm_group_bin_7281 (RW)
0x1ac: frame_vm_group_bin_0159 (RW)
0x1ad: frame_vm_group_bin_16310 (RW)
0x1ae: frame_vm_group_bin_9135 (RW)
0x1af: frame_vm_group_bin_1947 (RW)
0x1b0: frame_vm_group_bin_18045 (RW)
0x1b1: frame_vm_group_bin_10955 (RW)
0x1b2: frame_vm_group_bin_3770 (RW)
0x1b3: frame_vm_group_bin_19870 (RW)
0x1b4: frame_vm_group_bin_12684 (RW)
0x1b5: frame_vm_group_bin_5604 (RW)
0x1b6: frame_vm_group_bin_21702 (RW)
0x1b7: frame_vm_group_bin_14528 (RW)
0x1b8: frame_vm_group_bin_7313 (RW)
0x1b9: frame_vm_group_bin_0188 (RW)
0x1b: frame_vm_group_bin_7809 (RW)
0x1ba: frame_vm_group_bin_16343 (RW)
0x1bb: frame_vm_group_bin_9167 (RW)
0x1bc: frame_vm_group_bin_1980 (RW)
0x1bd: frame_vm_group_bin_18077 (RW)
0x1be: frame_vm_group_bin_10988 (RW)
0x1bf: frame_vm_group_bin_3803 (RW)
0x1c0: frame_vm_group_bin_19902 (RW)
0x1c1: frame_vm_group_bin_12712 (RW)
0x1c2: frame_vm_group_bin_5636 (RW)
0x1c3: frame_vm_group_bin_21736 (RW)
0x1c4: frame_vm_group_bin_14562 (RW)
0x1c5: frame_vm_group_bin_7347 (RW)
0x1c6: frame_vm_group_bin_0220 (RW)
0x1c7: frame_vm_group_bin_16376 (RW)
0x1c8: frame_vm_group_bin_9198 (RW)
0x1c9: frame_vm_group_bin_2013 (RW)
0x1c: frame_vm_group_bin_0954 (RW)
0x1ca: frame_vm_group_bin_18109 (RW)
0x1cb: frame_vm_group_bin_11021 (RW)
0x1cc: frame_vm_group_bin_3836 (RW)
0x1cd: frame_vm_group_bin_19934 (RW)
0x1ce: frame_vm_group_bin_12736 (RW)
0x1cf: frame_vm_group_bin_5669 (RW)
0x1d0: frame_vm_group_bin_21769 (RW)
0x1d1: frame_vm_group_bin_14595 (RW)
0x1d2: frame_vm_group_bin_7380 (RW)
0x1d3: frame_vm_group_bin_0245 (RW)
0x1d4: frame_vm_group_bin_16409 (RW)
0x1d5: frame_vm_group_bin_9223 (RW)
0x1d6: frame_vm_group_bin_2046 (RW)
0x1d7: frame_vm_group_bin_18142 (RW)
0x1d8: frame_vm_group_bin_11054 (RW)
0x1d9: frame_vm_group_bin_3869 (RW)
0x1d: frame_vm_group_bin_17148 (RW)
0x1da: frame_vm_group_bin_19968 (RW)
0x1db: frame_vm_group_bin_12767 (RW)
0x1dc: frame_vm_group_bin_5703 (RW)
0x1dd: frame_vm_group_bin_21803 (RW)
0x1de: frame_vm_group_bin_14628 (RW)
0x1df: frame_vm_group_bin_7414 (RW)
0x1e0: frame_vm_group_bin_0268 (RW)
0x1e1: frame_vm_group_bin_16443 (RW)
0x1e2: frame_vm_group_bin_9249 (RW)
0x1e3: frame_vm_group_bin_2080 (RW)
0x1e4: frame_vm_group_bin_18176 (RW)
0x1e5: frame_vm_group_bin_11088 (RW)
0x1e6: frame_vm_group_bin_3903 (RW)
0x1e7: frame_vm_group_bin_19999 (RW)
0x1e8: frame_vm_group_bin_12800 (RW)
0x1e9: frame_vm_group_bin_5735 (RW)
0x1e: frame_vm_group_bin_9938 (RW)
0x1ea: frame_vm_group_bin_21836 (RW)
0x1eb: frame_vm_group_bin_14661 (RW)
0x1ec: frame_vm_group_bin_7447 (RW)
0x1ed: frame_vm_group_bin_0295 (RW)
0x1ee: frame_vm_group_bin_16476 (RW)
0x1ef: frame_vm_group_bin_9271 (RW)
0x1f0: frame_vm_group_bin_2113 (RW)
0x1f1: frame_vm_group_bin_18208 (RW)
0x1f2: frame_vm_group_bin_11121 (RW)
0x1f3: frame_vm_group_bin_3936 (RW)
0x1f4: frame_vm_group_bin_20032 (RW)
0x1f5: frame_vm_group_bin_12832 (RW)
0x1f6: frame_vm_group_bin_5760 (RW)
0x1f7: frame_vm_group_bin_21869 (RW)
0x1f8: frame_vm_group_bin_14694 (RW)
0x1f9: frame_vm_group_bin_7480 (RW)
0x1f: frame_vm_group_bin_2780 (RW)
0x1fa: frame_vm_group_bin_0328 (RW)
0x1fb: frame_vm_group_bin_16510 (RW)
0x1fc: frame_vm_group_bin_9300 (RW)
0x1fd: frame_vm_group_bin_2148 (RW)
0x1fe: frame_vm_group_bin_18242 (RW)
0x1ff: frame_vm_group_bin_11154 (RW)
0x20: frame_vm_group_bin_18854 (RW)
0x21: frame_vm_group_bin_11734 (RW)
0x22: frame_vm_group_bin_4597 (RW)
0x23: frame_vm_group_bin_20706 (RW)
0x24: frame_vm_group_bin_13507 (RW)
0x25: frame_vm_group_bin_6321 (RW)
0x26: frame_vm_group_bin_22515 (RW)
0x27: frame_vm_group_bin_15332 (RW)
0x28: frame_vm_group_bin_8141 (RW)
0x29: frame_vm_group_bin_0987 (RW)
0x2: frame_vm_group_bin_0887 (RW)
0x2a: frame_vm_group_bin_17180 (RW)
0x2b: frame_vm_group_bin_9971 (RW)
0x2c: frame_vm_group_bin_2813 (RW)
0x2d: frame_vm_group_bin_18887 (RW)
0x2e: frame_vm_group_bin_11755 (RW)
0x2f: frame_vm_group_bin_4621 (RW)
0x30: frame_vm_group_bin_20739 (RW)
0x31: frame_vm_group_bin_13540 (RW)
0x32: frame_vm_group_bin_6354 (RW)
0x33: frame_vm_group_bin_22547 (RW)
0x34: frame_vm_group_bin_15365 (RW)
0x35: frame_vm_group_bin_8174 (RW)
0x36: frame_vm_group_bin_15747 (RW)
0x37: frame_vm_group_bin_17211 (RW)
0x38: frame_vm_group_bin_10004 (RW)
0x39: frame_vm_group_bin_2846 (RW)
0x3: frame_vm_group_bin_17082 (RW)
0x3a: frame_vm_group_bin_18921 (RW)
0x3b: frame_vm_group_bin_11781 (RW)
0x3c: frame_vm_group_bin_4652 (RW)
0x3d: frame_vm_group_bin_20773 (RW)
0x3e: frame_vm_group_bin_13574 (RW)
0x3f: frame_vm_group_bin_6385 (RW)
0x40: frame_vm_group_bin_22581 (RW)
0x41: frame_vm_group_bin_15399 (RW)
0x42: frame_vm_group_bin_8208 (RW)
0x43: frame_vm_group_bin_20390 (RW)
0x44: frame_vm_group_bin_17244 (RW)
0x45: frame_vm_group_bin_10038 (RW)
0x46: frame_vm_group_bin_2881 (RW)
0x47: frame_vm_group_bin_18953 (RW)
0x48: frame_vm_group_bin_11810 (RW)
0x49: frame_vm_group_bin_4684 (RW)
0x4: frame_vm_group_bin_9874 (RW)
0x4a: frame_vm_group_bin_20806 (RW)
0x4b: frame_vm_group_bin_13607 (RW)
0x4c: frame_vm_group_bin_6417 (RW)
0x4d: frame_vm_group_bin_22614 (RW)
0x4e: frame_vm_group_bin_15432 (RW)
0x4f: frame_vm_group_bin_8241 (RW)
0x50: frame_vm_group_bin_1062 (RW)
0x51: frame_vm_group_bin_17277 (RW)
0x52: frame_vm_group_bin_10071 (RW)
0x53: frame_vm_group_bin_2914 (RW)
0x54: frame_vm_group_bin_18984 (RW)
0x55: frame_vm_group_bin_11842 (RW)
0x56: frame_vm_group_bin_4716 (RW)
0x57: frame_vm_group_bin_20838 (RW)
0x58: frame_vm_group_bin_13639 (RW)
0x59: frame_vm_group_bin_6451 (RW)
0x5: frame_vm_group_bin_2713 (RW)
0x5a: frame_vm_group_bin_22648 (RW)
0x5b: frame_vm_group_bin_15466 (RW)
0x5c: frame_vm_group_bin_8274 (RW)
0x5d: frame_vm_group_bin_1090 (RW)
0x5e: frame_vm_group_bin_17311 (RW)
0x5f: frame_vm_group_bin_10105 (RW)
0x60: frame_vm_group_bin_2948 (RW)
0x61: frame_vm_group_bin_19018 (RW)
0x62: frame_vm_group_bin_11872 (RW)
0x63: frame_vm_group_bin_4749 (RW)
0x64: frame_vm_group_bin_20864 (RW)
0x65: frame_vm_group_bin_13673 (RW)
0x66: frame_vm_group_bin_6484 (RW)
0x67: frame_vm_group_bin_22681 (RW)
0x68: frame_vm_group_bin_15499 (RW)
0x69: frame_vm_group_bin_8307 (RW)
0x6: frame_vm_group_bin_18786 (RW)
0x6a: frame_vm_group_bin_1118 (RW)
0x6b: frame_vm_group_bin_17344 (RW)
0x6c: frame_vm_group_bin_10138 (RW)
0x6d: frame_vm_group_bin_2981 (RW)
0x6e: frame_vm_group_bin_19051 (RW)
0x6f: frame_vm_group_bin_11896 (RW)
0x70: frame_vm_group_bin_4782 (RW)
0x71: frame_vm_group_bin_20890 (RW)
0x72: frame_vm_group_bin_13706 (RW)
0x73: frame_vm_group_bin_6517 (RW)
0x74: frame_vm_group_bin_22714 (RW)
0x75: frame_vm_group_bin_15531 (RW)
0x76: frame_vm_group_bin_8340 (RW)
0x77: frame_vm_group_bin_1151 (RW)
0x78: frame_vm_group_bin_17376 (RW)
0x79: frame_vm_group_bin_10173 (RW)
0x7: frame_vm_group_bin_11681 (RW)
0x7a: frame_vm_group_bin_3015 (RW)
0x7b: frame_vm_group_bin_19085 (RW)
0x7c: frame_vm_group_bin_11923 (RW)
0x7d: frame_vm_group_bin_4815 (RW)
0x7e: frame_vm_group_bin_20919 (RW)
0x7f: frame_vm_group_bin_13739 (RW)
0x80: frame_vm_group_bin_6551 (RW)
0x81: frame_vm_group_bin_22747 (RW)
0x82: frame_vm_group_bin_15564 (RW)
0x83: frame_vm_group_bin_8374 (RW)
0x84: frame_vm_group_bin_1185 (RW)
0x85: frame_vm_group_bin_17405 (RW)
0x86: frame_vm_group_bin_10207 (RW)
0x87: frame_vm_group_bin_3048 (RW)
0x88: frame_vm_group_bin_19117 (RW)
0x89: frame_vm_group_bin_11953 (RW)
0x8: frame_vm_group_bin_4544 (RW)
0x8a: frame_vm_group_bin_4848 (RW)
0x8b: frame_vm_group_bin_20946 (RW)
0x8c: frame_vm_group_bin_13773 (RW)
0x8d: frame_vm_group_bin_6584 (RW)
0x8e: frame_vm_group_bin_22780 (RW)
0x8f: frame_vm_group_bin_15597 (RW)
0x90: frame_vm_group_bin_8407 (RW)
0x91: frame_vm_group_bin_1218 (RW)
0x92: frame_vm_group_bin_17429 (RW)
0x93: frame_vm_group_bin_10240 (RW)
0x94: frame_vm_group_bin_3081 (RW)
0x95: frame_vm_group_bin_19149 (RW)
0x96: frame_vm_group_bin_11986 (RW)
0x97: frame_vm_group_bin_4881 (RW)
0x98: frame_vm_group_bin_20974 (RW)
0x99: frame_vm_group_bin_13806 (RW)
0x9: frame_vm_group_bin_20640 (RW)
0x9a: frame_vm_group_bin_6618 (RW)
0x9b: frame_vm_group_bin_22814 (RW)
0x9c: frame_vm_group_bin_15631 (RW)
0x9d: frame_vm_group_bin_8441 (RW)
0x9e: frame_vm_group_bin_1251 (RW)
0x9f: frame_vm_group_bin_17457 (RW)
0xa0: frame_vm_group_bin_10274 (RW)
0xa1: frame_vm_group_bin_3114 (RW)
0xa2: frame_vm_group_bin_19183 (RW)
0xa3: frame_vm_group_bin_12018 (RW)
0xa4: frame_vm_group_bin_4915 (RW)
0xa5: frame_vm_group_bin_21008 (RW)
0xa6: frame_vm_group_bin_13836 (RW)
0xa7: frame_vm_group_bin_6651 (RW)
0xa8: frame_vm_group_bin_22847 (RW)
0xa9: frame_vm_group_bin_15664 (RW)
0xa: frame_vm_group_bin_13440 (RW)
0xaa: frame_vm_group_bin_8474 (RW)
0xab: frame_vm_group_bin_1282 (RW)
0xac: frame_vm_group_bin_17475 (RW)
0xad: frame_vm_group_bin_10307 (RW)
0xae: frame_vm_group_bin_3147 (RW)
0xaf: frame_vm_group_bin_19216 (RW)
0xb0: frame_vm_group_bin_12048 (RW)
0xb1: frame_vm_group_bin_4946 (RW)
0xb2: frame_vm_group_bin_21041 (RW)
0xb3: frame_vm_group_bin_13865 (RW)
0xb4: frame_vm_group_bin_6684 (RW)
0xb5: frame_vm_group_bin_22880 (RW)
0xb6: frame_vm_group_bin_15697 (RW)
0xb7: frame_vm_group_bin_8507 (RW)
0xb8: frame_vm_group_bin_1314 (RW)
0xb9: frame_vm_group_bin_17498 (RW)
0xb: frame_vm_group_bin_6256 (RW)
0xba: frame_vm_group_bin_10341 (RW)
0xbb: frame_vm_group_bin_3181 (RW)
0xbc: frame_vm_group_bin_19250 (RW)
0xbd: frame_vm_group_bin_12077 (RW)
0xbe: frame_vm_group_bin_4978 (RW)
0xbf: frame_vm_group_bin_21076 (RW)
0xc0: frame_vm_group_bin_13898 (RW)
0xc1: frame_vm_group_bin_6717 (RW)
0xc2: frame_vm_group_bin_22914 (RW)
0xc3: frame_vm_group_bin_15731 (RW)
0xc4: frame_vm_group_bin_8540 (RW)
0xc5: frame_vm_group_bin_1348 (RW)
0xc6: frame_vm_group_bin_17524 (RW)
0xc7: frame_vm_group_bin_10374 (RW)
0xc8: frame_vm_group_bin_3214 (RW)
0xc9: frame_vm_group_bin_19283 (RW)
0xc: frame_vm_group_bin_22448 (RW)
0xca: frame_vm_group_bin_12110 (RW)
0xcb: frame_vm_group_bin_5011 (RW)
0xcc: frame_vm_group_bin_21109 (RW)
0xcd: frame_vm_group_bin_13931 (RW)
0xce: frame_vm_group_bin_6750 (RW)
0xcf: frame_vm_group_bin_22947 (RW)
0xd0: frame_vm_group_bin_15764 (RW)
0xd1: frame_vm_group_bin_8571 (RW)
0xd2: frame_vm_group_bin_1382 (RW)
0xd3: frame_vm_group_bin_17549 (RW)
0xd4: frame_vm_group_bin_10401 (RW)
0xd5: frame_vm_group_bin_3246 (RW)
0xd6: frame_vm_group_bin_19316 (RW)
0xd7: frame_vm_group_bin_12142 (RW)
0xd8: frame_vm_group_bin_5044 (RW)
0xd9: frame_vm_group_bin_21141 (RW)
0xd: frame_vm_group_bin_15266 (RW)
0xda: frame_vm_group_bin_13965 (RW)
0xdb: frame_vm_group_bin_6783 (RW)
0xdc: frame_vm_group_bin_22980 (RW)
0xdd: frame_vm_group_bin_9318 (RW)
0xde: frame_vm_group_bin_8604 (RW)
0xdf: frame_vm_group_bin_1416 (RW)
0xe0: frame_vm_group_bin_17572 (RW)
0xe1: frame_vm_group_bin_10430 (RW)
0xe2: frame_vm_group_bin_3280 (RW)
0xe3: frame_vm_group_bin_19350 (RW)
0xe4: frame_vm_group_bin_12173 (RW)
0xe5: frame_vm_group_bin_5079 (RW)
0xe6: frame_vm_group_bin_21175 (RW)
0xe7: frame_vm_group_bin_13998 (RW)
0xe8: frame_vm_group_bin_16907 (RW)
0xe9: frame_vm_group_bin_23012 (RW)
0xe: frame_vm_group_bin_8076 (RW)
0xea: frame_vm_group_bin_15829 (RW)
0xeb: frame_vm_group_bin_8637 (RW)
0xec: frame_vm_group_bin_1449 (RW)
0xed: frame_vm_group_bin_17595 (RW)
0xee: frame_vm_group_bin_10460 (RW)
0xef: frame_vm_group_bin_3313 (RW)
0xf0: frame_vm_group_bin_19383 (RW)
0xf1: frame_vm_group_bin_12205 (RW)
0xf2: frame_vm_group_bin_5112 (RW)
0xf3: frame_vm_group_bin_21208 (RW)
0xf4: frame_vm_group_bin_14031 (RW)
0xf5: frame_vm_group_bin_6842 (RW)
0xf6: frame_vm_group_bin_23045 (RW)
0xf7: frame_vm_group_bin_15862 (RW)
0xf8: frame_vm_group_bin_8670 (RW)
0xf9: frame_vm_group_bin_1482 (RW)
0xf: frame_vm_group_bin_0920 (RW)
0xfa: frame_vm_group_bin_17623 (RW)
0xfb: frame_vm_group_bin_10494 (RW)
0xfc: frame_vm_group_bin_3347 (RW)
0xfd: frame_vm_group_bin_19416 (RW)
0xfe: frame_vm_group_bin_12235 (RW)
0xff: frame_vm_group_bin_5146 (RW)
}
pt_vm_group_bin_0044 {
0x0: frame_vm_group_bin_17749 (RW)
0x100: frame_vm_group_bin_0464 (RW)
0x101: frame_vm_group_bin_16654 (RW)
0x102: frame_vm_group_bin_9445 (RW)
0x103: frame_vm_group_bin_2285 (RW)
0x104: frame_vm_group_bin_18388 (RW)
0x105: frame_vm_group_bin_11300 (RW)
0x106: frame_vm_group_bin_4114 (RW)
0x107: frame_vm_group_bin_20209 (RW)
0x108: frame_vm_group_bin_13013 (RW)
0x109: frame_vm_group_bin_5888 (RW)
0x10: frame_vm_group_bin_19592 (RW)
0x10a: frame_vm_group_bin_22040 (RW)
0x10b: frame_vm_group_bin_14872 (RW)
0x10c: frame_vm_group_bin_7657 (RW)
0x10d: frame_vm_group_bin_0496 (RW)
0x10e: frame_vm_group_bin_16687 (RW)
0x10f: frame_vm_group_bin_9478 (RW)
0x110: frame_vm_group_bin_2318 (RW)
0x111: frame_vm_group_bin_18419 (RW)
0x112: frame_vm_group_bin_11333 (RW)
0x113: frame_vm_group_bin_4147 (RW)
0x114: frame_vm_group_bin_20242 (RW)
0x115: frame_vm_group_bin_13046 (RW)
0x116: frame_vm_group_bin_5914 (RW)
0x117: frame_vm_group_bin_7714 (RW)
0x118: frame_vm_group_bin_14905 (RW)
0x119: frame_vm_group_bin_7690 (RW)
0x11: frame_vm_group_bin_12412 (RW)
0x11a: frame_vm_group_bin_0529 (RW)
0x11b: frame_vm_group_bin_16721 (RW)
0x11c: frame_vm_group_bin_9512 (RW)
0x11d: frame_vm_group_bin_2352 (RW)
0x11e: frame_vm_group_bin_18453 (RW)
0x11f: frame_vm_group_bin_11365 (RW)
0x120: frame_vm_group_bin_4180 (RW)
0x121: frame_vm_group_bin_20275 (RW)
0x122: frame_vm_group_bin_13080 (RW)
0x123: frame_vm_group_bin_5938 (RW)
0x124: frame_vm_group_bin_12372 (RW)
0x125: frame_vm_group_bin_14939 (RW)
0x126: frame_vm_group_bin_7723 (RW)
0x127: frame_vm_group_bin_0560 (RW)
0x128: frame_vm_group_bin_16754 (RW)
0x129: frame_vm_group_bin_9545 (RW)
0x12: frame_vm_group_bin_5323 (RW)
0x12a: frame_vm_group_bin_2385 (RW)
0x12b: frame_vm_group_bin_18481 (RW)
0x12c: frame_vm_group_bin_11397 (RW)
0x12d: frame_vm_group_bin_4212 (RW)
0x12e: frame_vm_group_bin_20308 (RW)
0x12f: frame_vm_group_bin_13113 (RW)
0x130: frame_vm_group_bin_5963 (RW)
0x131: frame_vm_group_bin_22121 (RW)
0x132: frame_vm_group_bin_14972 (RW)
0x133: frame_vm_group_bin_7756 (RW)
0x134: frame_vm_group_bin_0592 (RW)
0x135: frame_vm_group_bin_16787 (RW)
0x136: frame_vm_group_bin_9578 (RW)
0x137: frame_vm_group_bin_2418 (RW)
0x138: frame_vm_group_bin_18508 (RW)
0x139: frame_vm_group_bin_11429 (RW)
0x13: frame_vm_group_bin_21418 (RW)
0x13a: frame_vm_group_bin_4246 (RW)
0x13b: frame_vm_group_bin_20344 (RW)
0x13c: frame_vm_group_bin_13147 (RW)
0x13d: frame_vm_group_bin_5992 (RW)
0x13e: frame_vm_group_bin_22155 (RW)
0x13f: frame_vm_group_bin_15006 (RW)
0x140: frame_vm_group_bin_7790 (RW)
0x141: frame_vm_group_bin_0624 (RW)
0x142: frame_vm_group_bin_16821 (RW)
0x143: frame_vm_group_bin_9612 (RW)
0x144: frame_vm_group_bin_2451 (RW)
0x145: frame_vm_group_bin_11711 (RW)
0x146: frame_vm_group_bin_11463 (RW)
0x147: frame_vm_group_bin_4279 (RW)
0x148: frame_vm_group_bin_20377 (RW)
0x149: frame_vm_group_bin_13180 (RW)
0x14: frame_vm_group_bin_14242 (RW)
0x14a: frame_vm_group_bin_6023 (RW)
0x14b: frame_vm_group_bin_22188 (RW)
0x14c: frame_vm_group_bin_15037 (RW)
0x14d: frame_vm_group_bin_7823 (RW)
0x14e: frame_vm_group_bin_0658 (RW)
0x14f: frame_vm_group_bin_16854 (RW)
0x150: frame_vm_group_bin_9645 (RW)
0x151: frame_vm_group_bin_2483 (RW)
0x152: frame_vm_group_bin_16389 (RW)
0x153: frame_vm_group_bin_11496 (RW)
0x154: frame_vm_group_bin_4312 (RW)
0x155: frame_vm_group_bin_20410 (RW)
0x156: frame_vm_group_bin_13213 (RW)
0x157: frame_vm_group_bin_6049 (RW)
0x158: frame_vm_group_bin_22221 (RW)
0x159: frame_vm_group_bin_6289 (RW)
0x15: frame_vm_group_bin_7029 (RW)
0x15a: frame_vm_group_bin_7856 (RW)
0x15b: frame_vm_group_bin_0692 (RW)
0x15c: frame_vm_group_bin_16887 (RW)
0x15d: frame_vm_group_bin_9679 (RW)
0x15e: frame_vm_group_bin_2517 (RW)
0x15f: frame_vm_group_bin_18594 (RW)
0x160: frame_vm_group_bin_11530 (RW)
0x161: frame_vm_group_bin_4348 (RW)
0x162: frame_vm_group_bin_20444 (RW)
0x163: frame_vm_group_bin_13247 (RW)
0x164: frame_vm_group_bin_6075 (RW)
0x165: frame_vm_group_bin_22255 (RW)
0x166: frame_vm_group_bin_11030 (RW)
0x167: frame_vm_group_bin_7889 (RW)
0x168: frame_vm_group_bin_0725 (RW)
0x169: frame_vm_group_bin_16919 (RW)
0x16: frame_vm_group_bin_3387 (RW)
0x16a: frame_vm_group_bin_9711 (RW)
0x16b: frame_vm_group_bin_2550 (RW)
0x16c: frame_vm_group_bin_18627 (RW)
0x16d: frame_vm_group_bin_11561 (RW)
0x16e: frame_vm_group_bin_4381 (RW)
0x16f: frame_vm_group_bin_20477 (RW)
0x170: frame_vm_group_bin_13280 (RW)
0x171: frame_vm_group_bin_6106 (RW)
0x172: frame_vm_group_bin_22287 (RW)
0x173: frame_vm_group_bin_15113 (RW)
0x174: frame_vm_group_bin_7922 (RW)
0x175: frame_vm_group_bin_0758 (RW)
0x176: frame_vm_group_bin_16952 (RW)
0x177: frame_vm_group_bin_9744 (RW)
0x178: frame_vm_group_bin_2583 (RW)
0x179: frame_vm_group_bin_18659 (RW)
0x17: frame_vm_group_bin_16076 (RW)
0x17a: frame_vm_group_bin_11589 (RW)
0x17b: frame_vm_group_bin_4415 (RW)
0x17c: frame_vm_group_bin_20511 (RW)
0x17d: frame_vm_group_bin_13314 (RW)
0x17e: frame_vm_group_bin_6139 (RW)
0x17f: frame_vm_group_bin_22321 (RW)
0x180: frame_vm_group_bin_20318 (RW)
0x181: frame_vm_group_bin_7957 (RW)
0x182: frame_vm_group_bin_0792 (RW)
0x183: frame_vm_group_bin_16986 (RW)
0x184: frame_vm_group_bin_9778 (RW)
0x185: frame_vm_group_bin_2617 (RW)
0x186: frame_vm_group_bin_18693 (RW)
0x187: frame_vm_group_bin_10316 (RW)
0x188: frame_vm_group_bin_4448 (RW)
0x189: frame_vm_group_bin_20544 (RW)
0x18: frame_vm_group_bin_8882 (RW)
0x18a: frame_vm_group_bin_13346 (RW)
0x18b: frame_vm_group_bin_6171 (RW)
0x18c: frame_vm_group_bin_22353 (RW)
0x18d: frame_vm_group_bin_15169 (RW)
0x18e: frame_vm_group_bin_7989 (RW)
0x18f: frame_vm_group_bin_0824 (RW)
0x190: frame_vm_group_bin_17019 (RW)
0x191: frame_vm_group_bin_9811 (RW)
0x192: frame_vm_group_bin_2650 (RW)
0x193: frame_vm_group_bin_18725 (RW)
0x194: frame_vm_group_bin_11636 (RW)
0x195: frame_vm_group_bin_4481 (RW)
0x196: frame_vm_group_bin_20577 (RW)
0x197: frame_vm_group_bin_13378 (RW)
0x198: frame_vm_group_bin_6202 (RW)
0x199: frame_vm_group_bin_22386 (RW)
0x19: frame_vm_group_bin_1694 (RW)
0x19a: frame_vm_group_bin_15203 (RW)
0x19b: frame_vm_group_bin_8020 (RW)
0x19c: frame_vm_group_bin_0858 (RW)
0x19d: frame_vm_group_bin_17053 (RW)
0x19e: frame_vm_group_bin_9845 (RW)
0x19f: frame_vm_group_bin_2684 (RW)
0x1: frame_vm_group_bin_10638 (RW)
0x1a0: frame_vm_group_bin_18757 (RW)
0x1a1: frame_vm_group_bin_19599 (RW)
0x1a2: frame_vm_group_bin_4515 (RW)
0x1a3: frame_vm_group_bin_20611 (RW)
0x1a4: frame_vm_group_bin_13411 (RW)
0x1a5: frame_vm_group_bin_6229 (RW)
0x1a6: frame_vm_group_bin_22419 (RW)
0x1a7: frame_vm_group_bin_15237 (RW)
0x1a8: frame_vm_group_bin_9582 (RW)
0x1a9: frame_vm_group_bin_0891 (RW)
0x1a: frame_vm_group_bin_20915 (RW)
0x1aa: frame_vm_group_bin_17086 (RW)
0x1ab: frame_vm_group_bin_9878 (RW)
0x1ac: frame_vm_group_bin_2717 (RW)
0x1ad: frame_vm_group_bin_18790 (RW)
0x1ae: frame_vm_group_bin_11683 (RW)
0x1af: frame_vm_group_bin_4548 (RW)
0x1b0: frame_vm_group_bin_20644 (RW)
0x1b1: frame_vm_group_bin_13444 (RW)
0x1b2: frame_vm_group_bin_6260 (RW)
0x1b3: frame_vm_group_bin_22452 (RW)
0x1b4: frame_vm_group_bin_15270 (RW)
0x1b5: frame_vm_group_bin_8080 (RW)
0x1b6: frame_vm_group_bin_0924 (RW)
0x1b7: frame_vm_group_bin_17119 (RW)
0x1b8: frame_vm_group_bin_9910 (RW)
0x1b9: frame_vm_group_bin_2750 (RW)
0x1b: frame_vm_group_bin_10703 (RW)
0x1ba: frame_vm_group_bin_18826 (RW)
0x1bb: frame_vm_group_bin_11712 (RW)
0x1bc: frame_vm_group_bin_4577 (RW)
0x1bd: frame_vm_group_bin_20677 (RW)
0x1be: frame_vm_group_bin_13478 (RW)
0x1bf: frame_vm_group_bin_6293 (RW)
0x1c0: frame_vm_group_bin_22486 (RW)
0x1c1: frame_vm_group_bin_15303 (RW)
0x1c2: frame_vm_group_bin_8112 (RW)
0x1c3: frame_vm_group_bin_0958 (RW)
0x1c4: frame_vm_group_bin_17152 (RW)
0x1c5: frame_vm_group_bin_9942 (RW)
0x1c6: frame_vm_group_bin_2784 (RW)
0x1c7: frame_vm_group_bin_18858 (RW)
0x1c8: frame_vm_group_bin_11736 (RW)
0x1c9: frame_vm_group_bin_8884 (RW)
0x1c: frame_vm_group_bin_3518 (RW)
0x1ca: frame_vm_group_bin_20710 (RW)
0x1cb: frame_vm_group_bin_13511 (RW)
0x1cc: frame_vm_group_bin_6325 (RW)
0x1cd: frame_vm_group_bin_22519 (RW)
0x1ce: frame_vm_group_bin_15336 (RW)
0x1cf: frame_vm_group_bin_8145 (RW)
0x1d0: frame_vm_group_bin_0991 (RW)
0x1d1: frame_vm_group_bin_17184 (RW)
0x1d2: frame_vm_group_bin_9975 (RW)
0x1d3: frame_vm_group_bin_2817 (RW)
0x1d4: frame_vm_group_bin_18891 (RW)
0x1d5: frame_vm_group_bin_11757 (RW)
0x1d6: frame_vm_group_bin_13522 (RW)
0x1d7: frame_vm_group_bin_20743 (RW)
0x1d8: frame_vm_group_bin_13544 (RW)
0x1d9: frame_vm_group_bin_6358 (RW)
0x1d: frame_vm_group_bin_19626 (RW)
0x1da: frame_vm_group_bin_22552 (RW)
0x1db: frame_vm_group_bin_15370 (RW)
0x1dc: frame_vm_group_bin_8179 (RW)
0x1dd: frame_vm_group_bin_1022 (RW)
0x1de: frame_vm_group_bin_17216 (RW)
0x1df: frame_vm_group_bin_10009 (RW)
0x1e0: frame_vm_group_bin_2851 (RW)
0x1e1: frame_vm_group_bin_18925 (RW)
0x1e2: frame_vm_group_bin_11783 (RW)
0x1e3: frame_vm_group_bin_4656 (RW)
0x1e4: frame_vm_group_bin_20777 (RW)
0x1e5: frame_vm_group_bin_13578 (RW)
0x1e6: frame_vm_group_bin_6389 (RW)
0x1e7: frame_vm_group_bin_22585 (RW)
0x1e8: frame_vm_group_bin_15403 (RW)
0x1e9: frame_vm_group_bin_8212 (RW)
0x1e: frame_vm_group_bin_12445 (RW)
0x1ea: frame_vm_group_bin_8152 (RW)
0x1eb: frame_vm_group_bin_17248 (RW)
0x1ec: frame_vm_group_bin_10042 (RW)
0x1ed: frame_vm_group_bin_2885 (RW)
0x1ee: frame_vm_group_bin_18957 (RW)
0x1ef: frame_vm_group_bin_11814 (RW)
0x1f0: frame_vm_group_bin_4688 (RW)
0x1f1: frame_vm_group_bin_20810 (RW)
0x1f2: frame_vm_group_bin_13611 (RW)
0x1f3: frame_vm_group_bin_6421 (RW)
0x1f4: frame_vm_group_bin_22618 (RW)
0x1f5: frame_vm_group_bin_15436 (RW)
0x1f6: frame_vm_group_bin_8245 (RW)
0x1f7: frame_vm_group_bin_12788 (RW)
0x1f8: frame_vm_group_bin_17281 (RW)
0x1f9: frame_vm_group_bin_10075 (RW)
0x1f: frame_vm_group_bin_5355 (RW)
0x1fa: frame_vm_group_bin_2919 (RW)
0x1fb: frame_vm_group_bin_18989 (RW)
0x1fc: frame_vm_group_bin_11845 (RW)
0x1fd: frame_vm_group_bin_4268 (RW)
0x1fe: frame_vm_group_bin_20843 (RW)
0x1ff: frame_vm_group_bin_13644 (RW)
0x20: frame_vm_group_bin_21451 (RW)
0x21: frame_vm_group_bin_14275 (RW)
0x22: frame_vm_group_bin_7061 (RW)
0x23: frame_vm_group_bin_2119 (RW)
0x24: frame_vm_group_bin_16109 (RW)
0x25: frame_vm_group_bin_8915 (RW)
0x26: frame_vm_group_bin_1727 (RW)
0x27: frame_vm_group_bin_17839 (RW)
0x28: frame_vm_group_bin_10735 (RW)
0x29: frame_vm_group_bin_3549 (RW)
0x2: frame_vm_group_bin_8719 (RW)
0x2a: frame_vm_group_bin_19656 (RW)
0x2b: frame_vm_group_bin_12477 (RW)
0x2c: frame_vm_group_bin_5387 (RW)
0x2d: frame_vm_group_bin_21483 (RW)
0x2e: frame_vm_group_bin_14306 (RW)
0x2f: frame_vm_group_bin_7093 (RW)
0x30: frame_vm_group_bin_0024 (RW)
0x31: frame_vm_group_bin_16140 (RW)
0x32: frame_vm_group_bin_8947 (RW)
0x33: frame_vm_group_bin_1759 (RW)
0x34: frame_vm_group_bin_17865 (RW)
0x35: frame_vm_group_bin_10768 (RW)
0x36: frame_vm_group_bin_3581 (RW)
0x37: frame_vm_group_bin_2655 (RW)
0x38: frame_vm_group_bin_12510 (RW)
0x39: frame_vm_group_bin_5420 (RW)
0x3: frame_vm_group_bin_19558 (RW)
0x3a: frame_vm_group_bin_21516 (RW)
0x3b: frame_vm_group_bin_14340 (RW)
0x3c: frame_vm_group_bin_7126 (RW)
0x3d: frame_vm_group_bin_0047 (RW)
0x3e: frame_vm_group_bin_16174 (RW)
0x3f: frame_vm_group_bin_8981 (RW)
0x40: frame_vm_group_bin_1793 (RW)
0x41: frame_vm_group_bin_17896 (RW)
0x42: frame_vm_group_bin_10801 (RW)
0x43: frame_vm_group_bin_3616 (RW)
0x44: frame_vm_group_bin_19716 (RW)
0x45: frame_vm_group_bin_12544 (RW)
0x46: frame_vm_group_bin_5453 (RW)
0x47: frame_vm_group_bin_21549 (RW)
0x48: frame_vm_group_bin_14373 (RW)
0x49: frame_vm_group_bin_7158 (RW)
0x4: frame_vm_group_bin_12379 (RW)
0x4a: frame_vm_group_bin_0072 (RW)
0x4b: frame_vm_group_bin_16205 (RW)
0x4c: frame_vm_group_bin_9014 (RW)
0x4d: frame_vm_group_bin_1826 (RW)
0x4e: frame_vm_group_bin_17928 (RW)
0x4f: frame_vm_group_bin_10834 (RW)
0x50: frame_vm_group_bin_3649 (RW)
0x51: frame_vm_group_bin_19749 (RW)
0x52: frame_vm_group_bin_12577 (RW)
0x53: frame_vm_group_bin_5485 (RW)
0x54: frame_vm_group_bin_21582 (RW)
0x55: frame_vm_group_bin_14406 (RW)
0x56: frame_vm_group_bin_7193 (RW)
0x57: frame_vm_group_bin_0098 (RW)
0x58: frame_vm_group_bin_16232 (RW)
0x59: frame_vm_group_bin_9047 (RW)
0x5: frame_vm_group_bin_5291 (RW)
0x5a: frame_vm_group_bin_1860 (RW)
0x5b: frame_vm_group_bin_17960 (RW)
0x5c: frame_vm_group_bin_10868 (RW)
0x5d: frame_vm_group_bin_3683 (RW)
0x5e: frame_vm_group_bin_19783 (RW)
0x5f: frame_vm_group_bin_12611 (RW)
0x60: frame_vm_group_bin_5518 (RW)
0x61: frame_vm_group_bin_21616 (RW)
0x62: frame_vm_group_bin_14440 (RW)
0x63: frame_vm_group_bin_7227 (RW)
0x64: frame_vm_group_bin_0123 (RW)
0x65: frame_vm_group_bin_6568 (RW)
0x66: frame_vm_group_bin_9081 (RW)
0x67: frame_vm_group_bin_1893 (RW)
0x68: frame_vm_group_bin_17991 (RW)
0x69: frame_vm_group_bin_10901 (RW)
0x6: frame_vm_group_bin_21385 (RW)
0x6a: frame_vm_group_bin_3716 (RW)
0x6b: frame_vm_group_bin_19816 (RW)
0x6c: frame_vm_group_bin_12643 (RW)
0x6d: frame_vm_group_bin_5551 (RW)
0x6e: frame_vm_group_bin_21649 (RW)
0x6f: frame_vm_group_bin_14473 (RW)
0x70: frame_vm_group_bin_7260 (RW)
0x71: frame_vm_group_bin_0144 (RW)
0x72: frame_vm_group_bin_11314 (RW)
0x73: frame_vm_group_bin_9114 (RW)
0x74: frame_vm_group_bin_1926 (RW)
0x75: frame_vm_group_bin_18024 (RW)
0x76: frame_vm_group_bin_10934 (RW)
0x77: frame_vm_group_bin_3749 (RW)
0x78: frame_vm_group_bin_19849 (RW)
0x79: frame_vm_group_bin_12670 (RW)
0x7: frame_vm_group_bin_14209 (RW)
0x7a: frame_vm_group_bin_5584 (RW)
0x7b: frame_vm_group_bin_21682 (RW)
0x7c: frame_vm_group_bin_14508 (RW)
0x7d: frame_vm_group_bin_7293 (RW)
0x7e: frame_vm_group_bin_0168 (RW)
0x7f: frame_vm_group_bin_16322 (RW)
0x80: frame_vm_group_bin_9147 (RW)
0x81: frame_vm_group_bin_1959 (RW)
0x82: frame_vm_group_bin_18057 (RW)
0x83: frame_vm_group_bin_10967 (RW)
0x84: frame_vm_group_bin_3782 (RW)
0x85: frame_vm_group_bin_19882 (RW)
0x86: frame_vm_group_bin_5899 (RW)
0x87: frame_vm_group_bin_5615 (RW)
0x88: frame_vm_group_bin_21715 (RW)
0x89: frame_vm_group_bin_14541 (RW)
0x8: frame_vm_group_bin_6996 (RW)
0x8a: frame_vm_group_bin_7326 (RW)
0x8b: frame_vm_group_bin_0200 (RW)
0x8c: frame_vm_group_bin_16355 (RW)
0x8d: frame_vm_group_bin_9179 (RW)
0x8e: frame_vm_group_bin_1992 (RW)
0x8f: frame_vm_group_bin_18089 (RW)
0x90: frame_vm_group_bin_11000 (RW)
0x91: frame_vm_group_bin_3815 (RW)
0x92: frame_vm_group_bin_19914 (RW)
0x93: frame_vm_group_bin_10585 (RW)
0x94: frame_vm_group_bin_5648 (RW)
0x95: frame_vm_group_bin_21748 (RW)
0x96: frame_vm_group_bin_14574 (RW)
0x97: frame_vm_group_bin_7359 (RW)
0x98: frame_vm_group_bin_0229 (RW)
0x99: frame_vm_group_bin_16388 (RW)
0x9: frame_vm_group_bin_23216 (RW)
0x9a: frame_vm_group_bin_9208 (RW)
0x9b: frame_vm_group_bin_2026 (RW)
0x9c: frame_vm_group_bin_18122 (RW)
0x9d: frame_vm_group_bin_11034 (RW)
0x9e: frame_vm_group_bin_3849 (RW)
0x9f: frame_vm_group_bin_19947 (RW)
0xa0: frame_vm_group_bin_15226 (RW)
0xa1: frame_vm_group_bin_5682 (RW)
0xa2: frame_vm_group_bin_21781 (RW)
0xa3: frame_vm_group_bin_14607 (RW)
0xa4: frame_vm_group_bin_7393 (RW)
0xa5: frame_vm_group_bin_0252 (RW)
0xa6: frame_vm_group_bin_16422 (RW)
0xa7: frame_vm_group_bin_5236 (RW)
0xa8: frame_vm_group_bin_2059 (RW)
0xa9: frame_vm_group_bin_18155 (RW)
0xa: frame_vm_group_bin_16043 (RW)
0xaa: frame_vm_group_bin_11067 (RW)
0xab: frame_vm_group_bin_3882 (RW)
0xac: frame_vm_group_bin_19980 (RW)
0xad: frame_vm_group_bin_12779 (RW)
0xae: frame_vm_group_bin_5715 (RW)
0xaf: frame_vm_group_bin_21815 (RW)
0xb0: frame_vm_group_bin_14640 (RW)
0xb1: frame_vm_group_bin_7426 (RW)
0xb2: frame_vm_group_bin_0276 (RW)
0xb3: frame_vm_group_bin_16455 (RW)
0xb4: frame_vm_group_bin_9866 (RW)
0xb5: frame_vm_group_bin_2092 (RW)
0xb6: frame_vm_group_bin_18188 (RW)
0xb7: frame_vm_group_bin_11100 (RW)
0xb8: frame_vm_group_bin_3915 (RW)
0xb9: frame_vm_group_bin_20011 (RW)
0xb: frame_vm_group_bin_8850 (RW)
0xba: frame_vm_group_bin_12813 (RW)
0xbb: frame_vm_group_bin_5746 (RW)
0xbc: frame_vm_group_bin_21849 (RW)
0xbd: frame_vm_group_bin_14674 (RW)
0xbe: frame_vm_group_bin_7460 (RW)
0xbf: frame_vm_group_bin_0307 (RW)
0xc0: frame_vm_group_bin_16489 (RW)
0xc1: frame_vm_group_bin_14529 (RW)
0xc2: frame_vm_group_bin_2127 (RW)
0xc3: frame_vm_group_bin_18221 (RW)
0xc4: frame_vm_group_bin_11133 (RW)
0xc5: frame_vm_group_bin_3948 (RW)
0xc6: frame_vm_group_bin_20045 (RW)
0xc7: frame_vm_group_bin_12845 (RW)
0xc8: frame_vm_group_bin_4532 (RW)
0xc9: frame_vm_group_bin_21882 (RW)
0xc: frame_vm_group_bin_1661 (RW)
0xca: frame_vm_group_bin_14707 (RW)
0xcb: frame_vm_group_bin_7493 (RW)
0xcc: frame_vm_group_bin_0339 (RW)
0xcd: frame_vm_group_bin_16522 (RW)
0xce: frame_vm_group_bin_9311 (RW)
0xcf: frame_vm_group_bin_2160 (RW)
0xd0: frame_vm_group_bin_18254 (RW)
0xd1: frame_vm_group_bin_11166 (RW)
0xd2: frame_vm_group_bin_3981 (RW)
0xd3: frame_vm_group_bin_20078 (RW)
0xd4: frame_vm_group_bin_12878 (RW)
0xd5: frame_vm_group_bin_9165 (RW)
0xd6: frame_vm_group_bin_21915 (RW)
0xd7: frame_vm_group_bin_14739 (RW)
0xd8: frame_vm_group_bin_7525 (RW)
0xd9: frame_vm_group_bin_0370 (RW)
0xd: frame_vm_group_bin_17779 (RW)
0xda: frame_vm_group_bin_16555 (RW)
0xdb: frame_vm_group_bin_9344 (RW)
0xdc: frame_vm_group_bin_2193 (RW)
0xdd: frame_vm_group_bin_18288 (RW)
0xde: frame_vm_group_bin_11200 (RW)
0xdf: frame_vm_group_bin_4015 (RW)
0xe0: frame_vm_group_bin_20111 (RW)
0xe1: frame_vm_group_bin_12912 (RW)
0xe2: frame_vm_group_bin_5813 (RW)
0xe3: frame_vm_group_bin_21948 (RW)
0xe4: frame_vm_group_bin_14773 (RW)
0xe5: frame_vm_group_bin_7557 (RW)
0xe6: frame_vm_group_bin_0401 (RW)
0xe7: frame_vm_group_bin_16588 (RW)
0xe8: frame_vm_group_bin_9377 (RW)
0xe9: frame_vm_group_bin_2223 (RW)
0xe: frame_vm_group_bin_10669 (RW)
0xea: frame_vm_group_bin_18321 (RW)
0xeb: frame_vm_group_bin_11233 (RW)
0xec: frame_vm_group_bin_4048 (RW)
0xed: frame_vm_group_bin_20144 (RW)
0xee: frame_vm_group_bin_12944 (RW)
0xef: frame_vm_group_bin_5838 (RW)
0xf0: frame_vm_group_bin_21981 (RW)
0xf1: frame_vm_group_bin_14805 (RW)
0xf2: frame_vm_group_bin_7590 (RW)
0xf3: frame_vm_group_bin_0430 (RW)
0xf4: frame_vm_group_bin_16620 (RW)
0xf5: frame_vm_group_bin_9411 (RW)
0xf6: frame_vm_group_bin_2251 (RW)
0xf7: frame_vm_group_bin_18354 (RW)
0xf8: frame_vm_group_bin_11266 (RW)
0xf9: frame_vm_group_bin_4081 (RW)
0xf: frame_vm_group_bin_13358 (RW)
0xfa: frame_vm_group_bin_20177 (RW)
0xfb: frame_vm_group_bin_12978 (RW)
0xfc: frame_vm_group_bin_23186 (RW)
0xfd: frame_vm_group_bin_22014 (RW)
0xfe: frame_vm_group_bin_14839 (RW)
0xff: frame_vm_group_bin_7624 (RW)
}
pt_vm_group_bin_0051 {
0x0: frame_vm_group_bin_19204 (RW)
0x100: frame_vm_group_bin_1935 (RW)
0x101: frame_vm_group_bin_18033 (RW)
0x102: frame_vm_group_bin_10943 (RW)
0x103: frame_vm_group_bin_3758 (RW)
0x104: frame_vm_group_bin_19858 (RW)
0x105: frame_vm_group_bin_10267 (RW)
0x106: frame_vm_group_bin_5592 (RW)
0x107: frame_vm_group_bin_21690 (RW)
0x108: frame_vm_group_bin_14516 (RW)
0x109: frame_vm_group_bin_7301 (RW)
0x10: frame_vm_group_bin_21063 (RW)
0x10a: frame_vm_group_bin_0176 (RW)
0x10b: frame_vm_group_bin_16330 (RW)
0x10c: frame_vm_group_bin_9155 (RW)
0x10d: frame_vm_group_bin_1967 (RW)
0x10e: frame_vm_group_bin_18065 (RW)
0x10f: frame_vm_group_bin_10975 (RW)
0x110: frame_vm_group_bin_3790 (RW)
0x111: frame_vm_group_bin_19890 (RW)
0x112: frame_vm_group_bin_14930 (RW)
0x113: frame_vm_group_bin_5623 (RW)
0x114: frame_vm_group_bin_21723 (RW)
0x115: frame_vm_group_bin_14549 (RW)
0x116: frame_vm_group_bin_7334 (RW)
0x117: frame_vm_group_bin_0208 (RW)
0x118: frame_vm_group_bin_16363 (RW)
0x119: frame_vm_group_bin_9186 (RW)
0x11: frame_vm_group_bin_13885 (RW)
0x11a: frame_vm_group_bin_2001 (RW)
0x11b: frame_vm_group_bin_18099 (RW)
0x11c: frame_vm_group_bin_11009 (RW)
0x11d: frame_vm_group_bin_3824 (RW)
0x11e: frame_vm_group_bin_19923 (RW)
0x11f: frame_vm_group_bin_12727 (RW)
0x120: frame_vm_group_bin_5657 (RW)
0x121: frame_vm_group_bin_21757 (RW)
0x122: frame_vm_group_bin_14583 (RW)
0x123: frame_vm_group_bin_7368 (RW)
0x124: frame_vm_group_bin_0236 (RW)
0x125: frame_vm_group_bin_16397 (RW)
0x126: frame_vm_group_bin_9216 (RW)
0x127: frame_vm_group_bin_2034 (RW)
0x128: frame_vm_group_bin_18130 (RW)
0x129: frame_vm_group_bin_11042 (RW)
0x12: frame_vm_group_bin_6705 (RW)
0x12a: frame_vm_group_bin_3857 (RW)
0x12b: frame_vm_group_bin_19955 (RW)
0x12c: frame_vm_group_bin_12754 (RW)
0x12d: frame_vm_group_bin_5690 (RW)
0x12e: frame_vm_group_bin_21789 (RW)
0x12f: frame_vm_group_bin_14615 (RW)
0x130: frame_vm_group_bin_7401 (RW)
0x131: frame_vm_group_bin_0257 (RW)
0x132: frame_vm_group_bin_16430 (RW)
0x133: frame_vm_group_bin_14199 (RW)
0x134: frame_vm_group_bin_2067 (RW)
0x135: frame_vm_group_bin_18163 (RW)
0x136: frame_vm_group_bin_11075 (RW)
0x137: frame_vm_group_bin_3890 (RW)
0x138: frame_vm_group_bin_19988 (RW)
0x139: frame_vm_group_bin_12787 (RW)
0x13: frame_vm_group_bin_22901 (RW)
0x13a: frame_vm_group_bin_5724 (RW)
0x13b: frame_vm_group_bin_21824 (RW)
0x13c: frame_vm_group_bin_14649 (RW)
0x13d: frame_vm_group_bin_7435 (RW)
0x13e: frame_vm_group_bin_0284 (RW)
0x13f: frame_vm_group_bin_16464 (RW)
0x140: frame_vm_group_bin_18825 (RW)
0x141: frame_vm_group_bin_2101 (RW)
0x142: frame_vm_group_bin_18196 (RW)
0x143: frame_vm_group_bin_11109 (RW)
0x144: frame_vm_group_bin_3924 (RW)
0x145: frame_vm_group_bin_20020 (RW)
0x146: frame_vm_group_bin_12820 (RW)
0x147: frame_vm_group_bin_5753 (RW)
0x148: frame_vm_group_bin_21857 (RW)
0x149: frame_vm_group_bin_14682 (RW)
0x14: frame_vm_group_bin_15718 (RW)
0x14a: frame_vm_group_bin_7468 (RW)
0x14b: frame_vm_group_bin_0315 (RW)
0x14c: frame_vm_group_bin_16497 (RW)
0x14d: frame_vm_group_bin_9289 (RW)
0x14e: frame_vm_group_bin_2135 (RW)
0x14f: frame_vm_group_bin_18229 (RW)
0x150: frame_vm_group_bin_11141 (RW)
0x151: frame_vm_group_bin_3956 (RW)
0x152: frame_vm_group_bin_20053 (RW)
0x153: frame_vm_group_bin_12853 (RW)
0x154: frame_vm_group_bin_13474 (RW)
0x155: frame_vm_group_bin_21890 (RW)
0x156: frame_vm_group_bin_14715 (RW)
0x157: frame_vm_group_bin_7501 (RW)
0x158: frame_vm_group_bin_0346 (RW)
0x159: frame_vm_group_bin_16530 (RW)
0x15: frame_vm_group_bin_8527 (RW)
0x15a: frame_vm_group_bin_9319 (RW)
0x15b: frame_vm_group_bin_2169 (RW)
0x15c: frame_vm_group_bin_18263 (RW)
0x15d: frame_vm_group_bin_11175 (RW)
0x15e: frame_vm_group_bin_3990 (RW)
0x15f: frame_vm_group_bin_20087 (RW)
0x160: frame_vm_group_bin_12887 (RW)
0x161: frame_vm_group_bin_18119 (RW)
0x162: frame_vm_group_bin_21923 (RW)
0x163: frame_vm_group_bin_14748 (RW)
0x164: frame_vm_group_bin_7533 (RW)
0x165: frame_vm_group_bin_0379 (RW)
0x166: frame_vm_group_bin_16563 (RW)
0x167: frame_vm_group_bin_9352 (RW)
0x168: frame_vm_group_bin_2201 (RW)
0x169: frame_vm_group_bin_18296 (RW)
0x16: frame_vm_group_bin_1335 (RW)
0x16a: frame_vm_group_bin_11208 (RW)
0x16b: frame_vm_group_bin_4023 (RW)
0x16c: frame_vm_group_bin_20119 (RW)
0x16d: frame_vm_group_bin_12920 (RW)
0x16e: frame_vm_group_bin_5818 (RW)
0x16f: frame_vm_group_bin_21956 (RW)
0x170: frame_vm_group_bin_14780 (RW)
0x171: frame_vm_group_bin_7565 (RW)
0x172: frame_vm_group_bin_0407 (RW)
0x173: frame_vm_group_bin_16596 (RW)
0x174: frame_vm_group_bin_9385 (RW)
0x175: frame_vm_group_bin_12743 (RW)
0x176: frame_vm_group_bin_18329 (RW)
0x177: frame_vm_group_bin_11241 (RW)
0x178: frame_vm_group_bin_4056 (RW)
0x179: frame_vm_group_bin_20152 (RW)
0x17: frame_vm_group_bin_17513 (RW)
0x17a: frame_vm_group_bin_12953 (RW)
0x17b: frame_vm_group_bin_5844 (RW)
0x17c: frame_vm_group_bin_21990 (RW)
0x17d: frame_vm_group_bin_14814 (RW)
0x17e: frame_vm_group_bin_7599 (RW)
0x17f: frame_vm_group_bin_0439 (RW)
0x180: frame_vm_group_bin_16629 (RW)
0x181: frame_vm_group_bin_9420 (RW)
0x182: frame_vm_group_bin_2260 (RW)
0x183: frame_vm_group_bin_18363 (RW)
0x184: frame_vm_group_bin_11275 (RW)
0x185: frame_vm_group_bin_4090 (RW)
0x186: frame_vm_group_bin_20184 (RW)
0x187: frame_vm_group_bin_12986 (RW)
0x188: frame_vm_group_bin_5869 (RW)
0x189: frame_vm_group_bin_22021 (RW)
0x18: frame_vm_group_bin_10361 (RW)
0x18a: frame_vm_group_bin_14847 (RW)
0x18b: frame_vm_group_bin_7632 (RW)
0x18c: frame_vm_group_bin_0472 (RW)
0x18d: frame_vm_group_bin_16662 (RW)
0x18e: frame_vm_group_bin_9453 (RW)
0x18f: frame_vm_group_bin_2293 (RW)
0x190: frame_vm_group_bin_18395 (RW)
0x191: frame_vm_group_bin_11308 (RW)
0x192: frame_vm_group_bin_4122 (RW)
0x193: frame_vm_group_bin_20217 (RW)
0x194: frame_vm_group_bin_13021 (RW)
0x195: frame_vm_group_bin_5894 (RW)
0x196: frame_vm_group_bin_12052 (RW)
0x197: frame_vm_group_bin_14880 (RW)
0x198: frame_vm_group_bin_7665 (RW)
0x199: frame_vm_group_bin_0504 (RW)
0x19: frame_vm_group_bin_3201 (RW)
0x19a: frame_vm_group_bin_16696 (RW)
0x19b: frame_vm_group_bin_9487 (RW)
0x19c: frame_vm_group_bin_2327 (RW)
0x19d: frame_vm_group_bin_18428 (RW)
0x19e: frame_vm_group_bin_0597 (RW)
0x19f: frame_vm_group_bin_22505 (RW)
0x1: frame_vm_group_bin_12037 (RW)
0x1a0: frame_vm_group_bin_20251 (RW)
0x1a1: frame_vm_group_bin_13055 (RW)
0x1a2: frame_vm_group_bin_5922 (RW)
0x1a3: frame_vm_group_bin_16792 (RW)
0x1a4: frame_vm_group_bin_14914 (RW)
0x1a5: frame_vm_group_bin_7699 (RW)
0x1a6: frame_vm_group_bin_0537 (RW)
0x1a7: frame_vm_group_bin_16729 (RW)
0x1a8: frame_vm_group_bin_9520 (RW)
0x1a9: frame_vm_group_bin_2360 (RW)
0x1a: frame_vm_group_bin_19271 (RW)
0x1aa: frame_vm_group_bin_18460 (RW)
0x1ab: frame_vm_group_bin_11373 (RW)
0x1ac: frame_vm_group_bin_4188 (RW)
0x1ad: frame_vm_group_bin_20283 (RW)
0x1ae: frame_vm_group_bin_13088 (RW)
0x1af: frame_vm_group_bin_5944 (RW)
0x1b0: frame_vm_group_bin_22096 (RW)
0x1b1: frame_vm_group_bin_14947 (RW)
0x1b2: frame_vm_group_bin_7731 (RW)
0x1b3: frame_vm_group_bin_0568 (RW)
0x1b4: frame_vm_group_bin_16762 (RW)
0x1b5: frame_vm_group_bin_9553 (RW)
0x1b6: frame_vm_group_bin_2393 (RW)
0x1b7: frame_vm_group_bin_18487 (RW)
0x1b8: frame_vm_group_bin_11405 (RW)
0x1b9: frame_vm_group_bin_4220 (RW)
0x1b: frame_vm_group_bin_12098 (RW)
0x1ba: frame_vm_group_bin_20319 (RW)
0x1bb: frame_vm_group_bin_13122 (RW)
0x1bc: frame_vm_group_bin_4245 (RW)
0x1bd: frame_vm_group_bin_22130 (RW)
0x1be: frame_vm_group_bin_14981 (RW)
0x1bf: frame_vm_group_bin_7765 (RW)
0x1c0: frame_vm_group_bin_0601 (RW)
0x1c1: frame_vm_group_bin_16796 (RW)
0x1c2: frame_vm_group_bin_9587 (RW)
0x1c3: frame_vm_group_bin_2426 (RW)
0x1c4: frame_vm_group_bin_16079 (RW)
0x1c5: frame_vm_group_bin_11438 (RW)
0x1c6: frame_vm_group_bin_4254 (RW)
0x1c7: frame_vm_group_bin_20352 (RW)
0x1c8: frame_vm_group_bin_13155 (RW)
0x1c9: frame_vm_group_bin_6000 (RW)
0x1c: frame_vm_group_bin_4999 (RW)
0x1ca: frame_vm_group_bin_22163 (RW)
0x1cb: frame_vm_group_bin_15014 (RW)
0x1cc: frame_vm_group_bin_7798 (RW)
0x1cd: frame_vm_group_bin_0632 (RW)
0x1ce: frame_vm_group_bin_16829 (RW)
0x1cf: frame_vm_group_bin_9620 (RW)
0x1d0: frame_vm_group_bin_2459 (RW)
0x1d1: frame_vm_group_bin_20722 (RW)
0x1d2: frame_vm_group_bin_11471 (RW)
0x1d3: frame_vm_group_bin_4287 (RW)
0x1d4: frame_vm_group_bin_20385 (RW)
0x1d5: frame_vm_group_bin_13188 (RW)
0x1d6: frame_vm_group_bin_6031 (RW)
0x1d7: frame_vm_group_bin_22196 (RW)
0x1d8: frame_vm_group_bin_15042 (RW)
0x1d9: frame_vm_group_bin_9243 (RW)
0x1d: frame_vm_group_bin_21097 (RW)
0x1da: frame_vm_group_bin_0667 (RW)
0x1db: frame_vm_group_bin_16863 (RW)
0x1dc: frame_vm_group_bin_9654 (RW)
0x1dd: frame_vm_group_bin_2492 (RW)
0x1de: frame_vm_group_bin_18569 (RW)
0x1df: frame_vm_group_bin_11505 (RW)
0x1e0: frame_vm_group_bin_4321 (RW)
0x1e1: frame_vm_group_bin_20419 (RW)
0x1e2: frame_vm_group_bin_13222 (RW)
0x1e3: frame_vm_group_bin_6057 (RW)
0x1e4: frame_vm_group_bin_22230 (RW)
0x1e5: frame_vm_group_bin_15344 (RW)
0x1e6: frame_vm_group_bin_7864 (RW)
0x1e7: frame_vm_group_bin_0700 (RW)
0x1e8: frame_vm_group_bin_16894 (RW)
0x1e9: frame_vm_group_bin_9686 (RW)
0x1e: frame_vm_group_bin_13919 (RW)
0x1ea: frame_vm_group_bin_2525 (RW)
0x1eb: frame_vm_group_bin_18602 (RW)
0x1ec: frame_vm_group_bin_11538 (RW)
0x1ed: frame_vm_group_bin_4356 (RW)
0x1ee: frame_vm_group_bin_20452 (RW)
0x1ef: frame_vm_group_bin_13255 (RW)
0x1f0: frame_vm_group_bin_6083 (RW)
0x1f1: frame_vm_group_bin_22263 (RW)
0x1f2: frame_vm_group_bin_19989 (RW)
0x1f3: frame_vm_group_bin_7897 (RW)
0x1f4: frame_vm_group_bin_0733 (RW)
0x1f5: frame_vm_group_bin_16927 (RW)
0x1f6: frame_vm_group_bin_9719 (RW)
0x1f7: frame_vm_group_bin_2558 (RW)
0x1f8: frame_vm_group_bin_18635 (RW)
0x1f9: frame_vm_group_bin_11568 (RW)
0x1f: frame_vm_group_bin_6738 (RW)
0x1fa: frame_vm_group_bin_4390 (RW)
0x1fb: frame_vm_group_bin_20486 (RW)
0x1fc: frame_vm_group_bin_13289 (RW)
0x1fd: frame_vm_group_bin_6114 (RW)
0x1fe: frame_vm_group_bin_22296 (RW)
0x1ff: frame_vm_group_bin_15122 (RW)
0x20: frame_vm_group_bin_22935 (RW)
0x21: frame_vm_group_bin_15752 (RW)
0x22: frame_vm_group_bin_8559 (RW)
0x23: frame_vm_group_bin_1370 (RW)
0x24: frame_vm_group_bin_17540 (RW)
0x25: frame_vm_group_bin_10394 (RW)
0x26: frame_vm_group_bin_3234 (RW)
0x27: frame_vm_group_bin_19304 (RW)
0x28: frame_vm_group_bin_12130 (RW)
0x29: frame_vm_group_bin_5032 (RW)
0x2: frame_vm_group_bin_4934 (RW)
0x2a: frame_vm_group_bin_21130 (RW)
0x2b: frame_vm_group_bin_13952 (RW)
0x2c: frame_vm_group_bin_6770 (RW)
0x2d: frame_vm_group_bin_22967 (RW)
0x2e: frame_vm_group_bin_15785 (RW)
0x2f: frame_vm_group_bin_8592 (RW)
0x30: frame_vm_group_bin_1403 (RW)
0x31: frame_vm_group_bin_17561 (RW)
0x32: frame_vm_group_bin_9816 (RW)
0x33: frame_vm_group_bin_3267 (RW)
0x34: frame_vm_group_bin_19337 (RW)
0x35: frame_vm_group_bin_12162 (RW)
0x36: frame_vm_group_bin_5065 (RW)
0x37: frame_vm_group_bin_21162 (RW)
0x38: frame_vm_group_bin_13985 (RW)
0x39: frame_vm_group_bin_6803 (RW)
0x3: frame_vm_group_bin_21029 (RW)
0x3a: frame_vm_group_bin_21657 (RW)
0x3b: frame_vm_group_bin_15818 (RW)
0x3c: frame_vm_group_bin_8625 (RW)
0x3d: frame_vm_group_bin_1437 (RW)
0x3e: frame_vm_group_bin_15935 (RW)
0x3f: frame_vm_group_bin_10448 (RW)
0x40: frame_vm_group_bin_3301 (RW)
0x41: frame_vm_group_bin_19371 (RW)
0x42: frame_vm_group_bin_12193 (RW)
0x43: frame_vm_group_bin_5100 (RW)
0x44: frame_vm_group_bin_21196 (RW)
0x45: frame_vm_group_bin_14019 (RW)
0x46: frame_vm_group_bin_6834 (RW)
0x47: frame_vm_group_bin_23033 (RW)
0x48: frame_vm_group_bin_15850 (RW)
0x49: frame_vm_group_bin_8658 (RW)
0x4: frame_vm_group_bin_13856 (RW)
0x4a: frame_vm_group_bin_1470 (RW)
0x4b: frame_vm_group_bin_17610 (RW)
0x4c: frame_vm_group_bin_10481 (RW)
0x4d: frame_vm_group_bin_3334 (RW)
0x4e: frame_vm_group_bin_19404 (RW)
0x4f: frame_vm_group_bin_12223 (RW)
0x50: frame_vm_group_bin_5133 (RW)
0x51: frame_vm_group_bin_21229 (RW)
0x52: frame_vm_group_bin_14052 (RW)
0x53: frame_vm_group_bin_9119 (RW)
0x54: frame_vm_group_bin_23066 (RW)
0x55: frame_vm_group_bin_15883 (RW)
0x56: frame_vm_group_bin_8692 (RW)
0x57: frame_vm_group_bin_1503 (RW)
0x58: frame_vm_group_bin_17643 (RW)
0x59: frame_vm_group_bin_10514 (RW)
0x5: frame_vm_group_bin_6672 (RW)
0x5a: frame_vm_group_bin_3368 (RW)
0x5b: frame_vm_group_bin_20934 (RW)
0x5c: frame_vm_group_bin_12256 (RW)
0x5d: frame_vm_group_bin_5167 (RW)
0x5e: frame_vm_group_bin_21263 (RW)
0x5f: frame_vm_group_bin_14086 (RW)
0x60: frame_vm_group_bin_13757 (RW)
0x61: frame_vm_group_bin_23100 (RW)
0x62: frame_vm_group_bin_15917 (RW)
0x63: frame_vm_group_bin_8726 (RW)
0x64: frame_vm_group_bin_1537 (RW)
0x65: frame_vm_group_bin_17677 (RW)
0x66: frame_vm_group_bin_10547 (RW)
0x67: frame_vm_group_bin_3398 (RW)
0x68: frame_vm_group_bin_19467 (RW)
0x69: frame_vm_group_bin_12289 (RW)
0x6: frame_vm_group_bin_22868 (RW)
0x6a: frame_vm_group_bin_5200 (RW)
0x6b: frame_vm_group_bin_21296 (RW)
0x6c: frame_vm_group_bin_14119 (RW)
0x6d: frame_vm_group_bin_18402 (RW)
0x6e: frame_vm_group_bin_23133 (RW)
0x6f: frame_vm_group_bin_15950 (RW)
0x70: frame_vm_group_bin_8759 (RW)
0x71: frame_vm_group_bin_1570 (RW)
0x72: frame_vm_group_bin_17703 (RW)
0x73: frame_vm_group_bin_10580 (RW)
0x74: frame_vm_group_bin_8390 (RW)
0x75: frame_vm_group_bin_19500 (RW)
0x76: frame_vm_group_bin_12322 (RW)
0x77: frame_vm_group_bin_5233 (RW)
0x78: frame_vm_group_bin_2680 (RW)
0x79: frame_vm_group_bin_14152 (RW)
0x7: frame_vm_group_bin_15685 (RW)
0x7a: frame_vm_group_bin_6941 (RW)
0x7b: frame_vm_group_bin_23166 (RW)
0x7c: frame_vm_group_bin_15986 (RW)
0x7d: frame_vm_group_bin_8793 (RW)
0x7e: frame_vm_group_bin_1604 (RW)
0x7f: frame_vm_group_bin_17731 (RW)
0x80: frame_vm_group_bin_10614 (RW)
0x81: frame_vm_group_bin_13026 (RW)
0x82: frame_vm_group_bin_19534 (RW)
0x83: frame_vm_group_bin_12355 (RW)
0x84: frame_vm_group_bin_5267 (RW)
0x85: frame_vm_group_bin_21361 (RW)
0x86: frame_vm_group_bin_14185 (RW)
0x87: frame_vm_group_bin_6972 (RW)
0x88: frame_vm_group_bin_23198 (RW)
0x89: frame_vm_group_bin_16019 (RW)
0x8: frame_vm_group_bin_8495 (RW)
0x8a: frame_vm_group_bin_8826 (RW)
0x8b: frame_vm_group_bin_1637 (RW)
0x8c: frame_vm_group_bin_17758 (RW)
0x8d: frame_vm_group_bin_10646 (RW)
0x8e: frame_vm_group_bin_3470 (RW)
0x8f: frame_vm_group_bin_19567 (RW)
0x90: frame_vm_group_bin_12388 (RW)
0x91: frame_vm_group_bin_5300 (RW)
0x92: frame_vm_group_bin_21394 (RW)
0x93: frame_vm_group_bin_14218 (RW)
0x94: frame_vm_group_bin_7005 (RW)
0x95: frame_vm_group_bin_7667 (RW)
0x96: frame_vm_group_bin_16052 (RW)
0x97: frame_vm_group_bin_8859 (RW)
0x98: frame_vm_group_bin_1670 (RW)
0x99: frame_vm_group_bin_17788 (RW)
0x9: frame_vm_group_bin_1303 (RW)
0x9a: frame_vm_group_bin_10679 (RW)
0x9b: frame_vm_group_bin_3497 (RW)
0x9c: frame_vm_group_bin_19602 (RW)
0x9d: frame_vm_group_bin_12422 (RW)
0x9e: frame_vm_group_bin_5332 (RW)
0x9f: frame_vm_group_bin_21427 (RW)
0xa0: frame_vm_group_bin_14251 (RW)
0xa1: frame_vm_group_bin_7038 (RW)
0xa2: frame_vm_group_bin_12325 (RW)
0xa3: frame_vm_group_bin_16085 (RW)
0xa4: frame_vm_group_bin_8891 (RW)
0xa5: frame_vm_group_bin_1703 (RW)
0xa6: frame_vm_group_bin_17818 (RW)
0xa7: frame_vm_group_bin_10711 (RW)
0xa8: frame_vm_group_bin_3525 (RW)
0xa9: frame_vm_group_bin_19634 (RW)
0xa: frame_vm_group_bin_17488 (RW)
0xaa: frame_vm_group_bin_12453 (RW)
0xab: frame_vm_group_bin_5363 (RW)
0xac: frame_vm_group_bin_21459 (RW)
0xad: frame_vm_group_bin_14283 (RW)
0xae: frame_vm_group_bin_7069 (RW)
0xaf: frame_vm_group_bin_17074 (RW)
0xb0: frame_vm_group_bin_16117 (RW)
0xb1: frame_vm_group_bin_8923 (RW)
0xb2: frame_vm_group_bin_1735 (RW)
0xb3: frame_vm_group_bin_17846 (RW)
0xb4: frame_vm_group_bin_10743 (RW)
0xb5: frame_vm_group_bin_3557 (RW)
0xb6: frame_vm_group_bin_19662 (RW)
0xb7: frame_vm_group_bin_12485 (RW)
0xb8: frame_vm_group_bin_5395 (RW)
0xb9: frame_vm_group_bin_21491 (RW)
0xb: frame_vm_group_bin_10328 (RW)
0xba: frame_vm_group_bin_14315 (RW)
0xbb: frame_vm_group_bin_7102 (RW)
0xbc: frame_vm_group_bin_0030 (RW)
0xbd: frame_vm_group_bin_16149 (RW)
0xbe: frame_vm_group_bin_8956 (RW)
0xbf: frame_vm_group_bin_1768 (RW)
0xc0: frame_vm_group_bin_17873 (RW)
0xc1: frame_vm_group_bin_10776 (RW)
0xc2: frame_vm_group_bin_3591 (RW)
0xc3: frame_vm_group_bin_19691 (RW)
0xc4: frame_vm_group_bin_12519 (RW)
0xc5: frame_vm_group_bin_5429 (RW)
0xc6: frame_vm_group_bin_21524 (RW)
0xc7: frame_vm_group_bin_14348 (RW)
0xc8: frame_vm_group_bin_7133 (RW)
0xc9: frame_vm_group_bin_0053 (RW)
0xc: frame_vm_group_bin_3168 (RW)
0xca: frame_vm_group_bin_16182 (RW)
0xcb: frame_vm_group_bin_8989 (RW)
0xcc: frame_vm_group_bin_1801 (RW)
0xcd: frame_vm_group_bin_17904 (RW)
0xce: frame_vm_group_bin_10809 (RW)
0xcf: frame_vm_group_bin_3624 (RW)
0xd0: frame_vm_group_bin_19724 (RW)
0xd1: frame_vm_group_bin_12552 (RW)
0xd2: frame_vm_group_bin_5461 (RW)
0xd3: frame_vm_group_bin_21557 (RW)
0xd4: frame_vm_group_bin_14381 (RW)
0xd5: frame_vm_group_bin_7166 (RW)
0xd6: frame_vm_group_bin_0079 (RW)
0xd7: frame_vm_group_bin_16212 (RW)
0xd8: frame_vm_group_bin_9022 (RW)
0xd9: frame_vm_group_bin_1834 (RW)
0xd: frame_vm_group_bin_19237 (RW)
0xda: frame_vm_group_bin_17936 (RW)
0xdb: frame_vm_group_bin_10843 (RW)
0xdc: frame_vm_group_bin_3658 (RW)
0xdd: frame_vm_group_bin_19758 (RW)
0xde: frame_vm_group_bin_12586 (RW)
0xdf: frame_vm_group_bin_5494 (RW)
0xe0: frame_vm_group_bin_21591 (RW)
0xe1: frame_vm_group_bin_14415 (RW)
0xe2: frame_vm_group_bin_7202 (RW)
0xe3: frame_vm_group_bin_0105 (RW)
0xe4: frame_vm_group_bin_10983 (RW)
0xe5: frame_vm_group_bin_9056 (RW)
0xe6: frame_vm_group_bin_1868 (RW)
0xe7: frame_vm_group_bin_17968 (RW)
0xe8: frame_vm_group_bin_10875 (RW)
0xe9: frame_vm_group_bin_3691 (RW)
0xe: frame_vm_group_bin_12064 (RW)
0xea: frame_vm_group_bin_19791 (RW)
0xeb: frame_vm_group_bin_12619 (RW)
0xec: frame_vm_group_bin_5526 (RW)
0xed: frame_vm_group_bin_21624 (RW)
0xee: frame_vm_group_bin_14448 (RW)
0xef: frame_vm_group_bin_7235 (RW)
0xf0: frame_vm_group_bin_0128 (RW)
0xf1: frame_vm_group_bin_15628 (RW)
0xf2: frame_vm_group_bin_9089 (RW)
0xf3: frame_vm_group_bin_1901 (RW)
0xf4: frame_vm_group_bin_17999 (RW)
0xf5: frame_vm_group_bin_10909 (RW)
0xf6: frame_vm_group_bin_3724 (RW)
0xf7: frame_vm_group_bin_19824 (RW)
0xf8: frame_vm_group_bin_12650 (RW)
0xf9: frame_vm_group_bin_5559 (RW)
0xf: frame_vm_group_bin_4965 (RW)
0xfa: frame_vm_group_bin_21658 (RW)
0xfb: frame_vm_group_bin_14482 (RW)
0xfc: frame_vm_group_bin_7269 (RW)
0xfd: frame_vm_group_bin_0150 (RW)
0xfe: frame_vm_group_bin_16298 (RW)
0xff: frame_vm_group_bin_9123 (RW)
}
pt_vm_group_bin_0054 {
0x0: frame_vm_group_bin_11629 (RW)
0x100: frame_vm_group_bin_17588 (RW)
0x101: frame_vm_group_bin_10450 (RW)
0x102: frame_vm_group_bin_3303 (RW)
0x103: frame_vm_group_bin_19373 (RW)
0x104: frame_vm_group_bin_12195 (RW)
0x105: frame_vm_group_bin_5102 (RW)
0x106: frame_vm_group_bin_21198 (RW)
0x107: frame_vm_group_bin_14021 (RW)
0x108: frame_vm_group_bin_17584 (RW)
0x109: frame_vm_group_bin_23035 (RW)
0x10: frame_vm_group_bin_13396 (RW)
0x10a: frame_vm_group_bin_15852 (RW)
0x10b: frame_vm_group_bin_8660 (RW)
0x10c: frame_vm_group_bin_1472 (RW)
0x10d: frame_vm_group_bin_17612 (RW)
0x10e: frame_vm_group_bin_10483 (RW)
0x10f: frame_vm_group_bin_3336 (RW)
0x110: frame_vm_group_bin_19406 (RW)
0x111: frame_vm_group_bin_12225 (RW)
0x112: frame_vm_group_bin_5135 (RW)
0x113: frame_vm_group_bin_21231 (RW)
0x114: frame_vm_group_bin_14054 (RW)
0x115: frame_vm_group_bin_6861 (RW)
0x116: frame_vm_group_bin_23068 (RW)
0x117: frame_vm_group_bin_15885 (RW)
0x118: frame_vm_group_bin_8694 (RW)
0x119: frame_vm_group_bin_1505 (RW)
0x11: frame_vm_group_bin_6216 (RW)
0x11a: frame_vm_group_bin_17646 (RW)
0x11b: frame_vm_group_bin_13640 (RW)
0x11c: frame_vm_group_bin_3370 (RW)
0x11d: frame_vm_group_bin_19437 (RW)
0x11e: frame_vm_group_bin_12258 (RW)
0x11f: frame_vm_group_bin_5169 (RW)
0x120: frame_vm_group_bin_21265 (RW)
0x121: frame_vm_group_bin_14088 (RW)
0x122: frame_vm_group_bin_6887 (RW)
0x123: frame_vm_group_bin_23102 (RW)
0x124: frame_vm_group_bin_15919 (RW)
0x125: frame_vm_group_bin_8728 (RW)
0x126: frame_vm_group_bin_1539 (RW)
0x127: frame_vm_group_bin_17679 (RW)
0x128: frame_vm_group_bin_10549 (RW)
0x129: frame_vm_group_bin_16932 (RW)
0x12: frame_vm_group_bin_22405 (RW)
0x12a: frame_vm_group_bin_19469 (RW)
0x12b: frame_vm_group_bin_12291 (RW)
0x12c: frame_vm_group_bin_5202 (RW)
0x12d: frame_vm_group_bin_21298 (RW)
0x12e: frame_vm_group_bin_14121 (RW)
0x12f: frame_vm_group_bin_6911 (RW)
0x130: frame_vm_group_bin_23135 (RW)
0x131: frame_vm_group_bin_15952 (RW)
0x132: frame_vm_group_bin_8761 (RW)
0x133: frame_vm_group_bin_1572 (RW)
0x134: frame_vm_group_bin_17705 (RW)
0x135: frame_vm_group_bin_10582 (RW)
0x136: frame_vm_group_bin_3422 (RW)
0x137: frame_vm_group_bin_19502 (RW)
0x138: frame_vm_group_bin_18637 (RW)
0x139: frame_vm_group_bin_5235 (RW)
0x13: frame_vm_group_bin_15221 (RW)
0x13a: frame_vm_group_bin_21330 (RW)
0x13b: frame_vm_group_bin_14155 (RW)
0x13c: frame_vm_group_bin_6943 (RW)
0x13d: frame_vm_group_bin_23168 (RW)
0x13e: frame_vm_group_bin_15988 (RW)
0x13f: frame_vm_group_bin_8795 (RW)
0x140: frame_vm_group_bin_1606 (RW)
0x141: frame_vm_group_bin_17733 (RW)
0x142: frame_vm_group_bin_10616 (RW)
0x143: frame_vm_group_bin_3445 (RW)
0x144: frame_vm_group_bin_19536 (RW)
0x145: frame_vm_group_bin_12357 (RW)
0x146: frame_vm_group_bin_5269 (RW)
0x147: frame_vm_group_bin_21363 (RW)
0x148: frame_vm_group_bin_14187 (RW)
0x149: frame_vm_group_bin_6974 (RW)
0x14: frame_vm_group_bin_8034 (RW)
0x14a: frame_vm_group_bin_23200 (RW)
0x14b: frame_vm_group_bin_16021 (RW)
0x14c: frame_vm_group_bin_8828 (RW)
0x14d: frame_vm_group_bin_1639 (RW)
0x14e: frame_vm_group_bin_17760 (RW)
0x14f: frame_vm_group_bin_10648 (RW)
0x150: frame_vm_group_bin_3471 (RW)
0x151: frame_vm_group_bin_19569 (RW)
0x152: frame_vm_group_bin_12390 (RW)
0x153: frame_vm_group_bin_5302 (RW)
0x154: frame_vm_group_bin_21396 (RW)
0x155: frame_vm_group_bin_14220 (RW)
0x156: frame_vm_group_bin_7007 (RW)
0x157: frame_vm_group_bin_20859 (RW)
0x158: frame_vm_group_bin_16054 (RW)
0x159: frame_vm_group_bin_17935 (RW)
0x15: frame_vm_group_bin_0876 (RW)
0x15a: frame_vm_group_bin_1673 (RW)
0x15b: frame_vm_group_bin_17790 (RW)
0x15c: frame_vm_group_bin_10681 (RW)
0x15d: frame_vm_group_bin_3499 (RW)
0x15e: frame_vm_group_bin_19604 (RW)
0x15f: frame_vm_group_bin_12424 (RW)
0x160: frame_vm_group_bin_5334 (RW)
0x161: frame_vm_group_bin_21429 (RW)
0x162: frame_vm_group_bin_14253 (RW)
0x163: frame_vm_group_bin_7040 (RW)
0x164: frame_vm_group_bin_23244 (RW)
0x165: frame_vm_group_bin_16087 (RW)
0x166: frame_vm_group_bin_8893 (RW)
0x167: frame_vm_group_bin_1705 (RW)
0x168: frame_vm_group_bin_17820 (RW)
0x169: frame_vm_group_bin_10713 (RW)
0x16: frame_vm_group_bin_17071 (RW)
0x16a: frame_vm_group_bin_3527 (RW)
0x16b: frame_vm_group_bin_19636 (RW)
0x16c: frame_vm_group_bin_12455 (RW)
0x16d: frame_vm_group_bin_5365 (RW)
0x16e: frame_vm_group_bin_21461 (RW)
0x16f: frame_vm_group_bin_14285 (RW)
0x170: frame_vm_group_bin_7071 (RW)
0x171: frame_vm_group_bin_6844 (RW)
0x172: frame_vm_group_bin_16119 (RW)
0x173: frame_vm_group_bin_8925 (RW)
0x174: frame_vm_group_bin_1737 (RW)
0x175: frame_vm_group_bin_17848 (RW)
0x176: frame_vm_group_bin_10745 (RW)
0x177: frame_vm_group_bin_3559 (RW)
0x178: frame_vm_group_bin_17451 (RW)
0x179: frame_vm_group_bin_12487 (RW)
0x17: frame_vm_group_bin_9863 (RW)
0x17a: frame_vm_group_bin_5398 (RW)
0x17b: frame_vm_group_bin_15863 (RW)
0x17c: frame_vm_group_bin_14317 (RW)
0x17d: frame_vm_group_bin_7104 (RW)
0x17e: frame_vm_group_bin_0032 (RW)
0x17f: frame_vm_group_bin_16151 (RW)
0x180: frame_vm_group_bin_8958 (RW)
0x181: frame_vm_group_bin_1770 (RW)
0x182: frame_vm_group_bin_17875 (RW)
0x183: frame_vm_group_bin_10778 (RW)
0x184: frame_vm_group_bin_3593 (RW)
0x185: frame_vm_group_bin_19693 (RW)
0x186: frame_vm_group_bin_12521 (RW)
0x187: frame_vm_group_bin_5431 (RW)
0x188: frame_vm_group_bin_21526 (RW)
0x189: frame_vm_group_bin_14350 (RW)
0x18: frame_vm_group_bin_2702 (RW)
0x18a: frame_vm_group_bin_7135 (RW)
0x18b: frame_vm_group_bin_0055 (RW)
0x18c: frame_vm_group_bin_16184 (RW)
0x18d: frame_vm_group_bin_8991 (RW)
0x18e: frame_vm_group_bin_1803 (RW)
0x18f: frame_vm_group_bin_17906 (RW)
0x190: frame_vm_group_bin_10811 (RW)
0x191: frame_vm_group_bin_3626 (RW)
0x192: frame_vm_group_bin_19726 (RW)
0x193: frame_vm_group_bin_12554 (RW)
0x194: frame_vm_group_bin_5463 (RW)
0x195: frame_vm_group_bin_21559 (RW)
0x196: frame_vm_group_bin_14383 (RW)
0x197: frame_vm_group_bin_7168 (RW)
0x198: frame_vm_group_bin_0081 (RW)
0x199: frame_vm_group_bin_16214 (RW)
0x19: frame_vm_group_bin_18775 (RW)
0x19a: frame_vm_group_bin_9025 (RW)
0x19b: frame_vm_group_bin_1837 (RW)
0x19c: frame_vm_group_bin_17938 (RW)
0x19d: frame_vm_group_bin_10845 (RW)
0x19e: frame_vm_group_bin_3660 (RW)
0x19f: frame_vm_group_bin_19760 (RW)
0x1: frame_vm_group_bin_4467 (RW)
0x1a0: frame_vm_group_bin_12588 (RW)
0x1a1: frame_vm_group_bin_5496 (RW)
0x1a2: frame_vm_group_bin_21593 (RW)
0x1a3: frame_vm_group_bin_14417 (RW)
0x1a4: frame_vm_group_bin_7204 (RW)
0x1a5: frame_vm_group_bin_0107 (RW)
0x1a6: frame_vm_group_bin_16241 (RW)
0x1a7: frame_vm_group_bin_9058 (RW)
0x1a8: frame_vm_group_bin_1870 (RW)
0x1a9: frame_vm_group_bin_17970 (RW)
0x1a: frame_vm_group_bin_11672 (RW)
0x1aa: frame_vm_group_bin_10877 (RW)
0x1ab: frame_vm_group_bin_3693 (RW)
0x1ac: frame_vm_group_bin_19793 (RW)
0x1ad: frame_vm_group_bin_12621 (RW)
0x1ae: frame_vm_group_bin_5528 (RW)
0x1af: frame_vm_group_bin_21626 (RW)
0x1b0: frame_vm_group_bin_14450 (RW)
0x1b1: frame_vm_group_bin_7237 (RW)
0x1b2: frame_vm_group_bin_0130 (RW)
0x1b3: frame_vm_group_bin_16268 (RW)
0x1b4: frame_vm_group_bin_9091 (RW)
0x1b5: frame_vm_group_bin_1903 (RW)
0x1b6: frame_vm_group_bin_18001 (RW)
0x1b7: frame_vm_group_bin_10911 (RW)
0x1b8: frame_vm_group_bin_3726 (RW)
0x1b9: frame_vm_group_bin_19826 (RW)
0x1b: frame_vm_group_bin_4534 (RW)
0x1ba: frame_vm_group_bin_12653 (RW)
0x1bb: frame_vm_group_bin_5562 (RW)
0x1bc: frame_vm_group_bin_21660 (RW)
0x1bd: frame_vm_group_bin_14484 (RW)
0x1be: frame_vm_group_bin_7271 (RW)
0x1bf: frame_vm_group_bin_0152 (RW)
0x1c0: frame_vm_group_bin_16300 (RW)
0x1c1: frame_vm_group_bin_9125 (RW)
0x1c2: frame_vm_group_bin_1937 (RW)
0x1c3: frame_vm_group_bin_18035 (RW)
0x1c4: frame_vm_group_bin_10945 (RW)
0x1c5: frame_vm_group_bin_3760 (RW)
0x1c6: frame_vm_group_bin_19860 (RW)
0x1c7: frame_vm_group_bin_0118 (RW)
0x1c8: frame_vm_group_bin_5594 (RW)
0x1c9: frame_vm_group_bin_21692 (RW)
0x1c: frame_vm_group_bin_20630 (RW)
0x1ca: frame_vm_group_bin_14518 (RW)
0x1cb: frame_vm_group_bin_7303 (RW)
0x1cc: frame_vm_group_bin_0178 (RW)
0x1cd: frame_vm_group_bin_16332 (RW)
0x1ce: frame_vm_group_bin_9157 (RW)
0x1cf: frame_vm_group_bin_1969 (RW)
0x1d0: frame_vm_group_bin_18067 (RW)
0x1d1: frame_vm_group_bin_10977 (RW)
0x1d2: frame_vm_group_bin_3792 (RW)
0x1d3: frame_vm_group_bin_19892 (RW)
0x1d4: frame_vm_group_bin_12701 (RW)
0x1d5: frame_vm_group_bin_5625 (RW)
0x1d6: frame_vm_group_bin_21725 (RW)
0x1d7: frame_vm_group_bin_14551 (RW)
0x1d8: frame_vm_group_bin_7336 (RW)
0x1d9: frame_vm_group_bin_0210 (RW)
0x1d: frame_vm_group_bin_13430 (RW)
0x1da: frame_vm_group_bin_16366 (RW)
0x1db: frame_vm_group_bin_9189 (RW)
0x1dc: frame_vm_group_bin_2003 (RW)
0x1dd: frame_vm_group_bin_18100 (RW)
0x1de: frame_vm_group_bin_11011 (RW)
0x1df: frame_vm_group_bin_3826 (RW)
0x1e0: frame_vm_group_bin_19924 (RW)
0x1e1: frame_vm_group_bin_12728 (RW)
0x1e2: frame_vm_group_bin_5659 (RW)
0x1e3: frame_vm_group_bin_21759 (RW)
0x1e4: frame_vm_group_bin_14585 (RW)
0x1e5: frame_vm_group_bin_7370 (RW)
0x1e6: frame_vm_group_bin_0238 (RW)
0x1e7: frame_vm_group_bin_16399 (RW)
0x1e8: frame_vm_group_bin_22717 (RW)
0x1e9: frame_vm_group_bin_2036 (RW)
0x1e: frame_vm_group_bin_6246 (RW)
0x1ea: frame_vm_group_bin_18132 (RW)
0x1eb: frame_vm_group_bin_11044 (RW)
0x1ec: frame_vm_group_bin_3859 (RW)
0x1ed: frame_vm_group_bin_19957 (RW)
0x1ee: frame_vm_group_bin_12756 (RW)
0x1ef: frame_vm_group_bin_5692 (RW)
0x1f0: frame_vm_group_bin_21791 (RW)
0x1f1: frame_vm_group_bin_14617 (RW)
0x1f2: frame_vm_group_bin_7403 (RW)
0x1f3: frame_vm_group_bin_0259 (RW)
0x1f4: frame_vm_group_bin_16432 (RW)
0x1f5: frame_vm_group_bin_9240 (RW)
0x1f6: frame_vm_group_bin_2069 (RW)
0x1f7: frame_vm_group_bin_18165 (RW)
0x1f8: frame_vm_group_bin_11077 (RW)
0x1f9: frame_vm_group_bin_3892 (RW)
0x1f: frame_vm_group_bin_22438 (RW)
0x1fa: frame_vm_group_bin_19990 (RW)
0x1fb: frame_vm_group_bin_12790 (RW)
0x1fc: frame_vm_group_bin_5726 (RW)
0x1fd: frame_vm_group_bin_21826 (RW)
0x1fe: frame_vm_group_bin_14651 (RW)
0x1ff: frame_vm_group_bin_7437 (RW)
0x20: frame_vm_group_bin_15256 (RW)
0x21: frame_vm_group_bin_8066 (RW)
0x22: frame_vm_group_bin_0910 (RW)
0x23: frame_vm_group_bin_17105 (RW)
0x24: frame_vm_group_bin_9896 (RW)
0x25: frame_vm_group_bin_2736 (RW)
0x26: frame_vm_group_bin_18809 (RW)
0x27: frame_vm_group_bin_11699 (RW)
0x28: frame_vm_group_bin_4566 (RW)
0x29: frame_vm_group_bin_20662 (RW)
0x2: frame_vm_group_bin_20563 (RW)
0x2a: frame_vm_group_bin_13463 (RW)
0x2b: frame_vm_group_bin_6278 (RW)
0x2c: frame_vm_group_bin_22471 (RW)
0x2d: frame_vm_group_bin_15288 (RW)
0x2e: frame_vm_group_bin_8098 (RW)
0x2f: frame_vm_group_bin_0943 (RW)
0x30: frame_vm_group_bin_17138 (RW)
0x31: frame_vm_group_bin_9929 (RW)
0x32: frame_vm_group_bin_2769 (RW)
0x33: frame_vm_group_bin_18843 (RW)
0x34: frame_vm_group_bin_11726 (RW)
0x35: frame_vm_group_bin_17212 (RW)
0x36: frame_vm_group_bin_20695 (RW)
0x37: frame_vm_group_bin_13496 (RW)
0x38: frame_vm_group_bin_6311 (RW)
0x39: frame_vm_group_bin_22504 (RW)
0x3: frame_vm_group_bin_13365 (RW)
0x3a: frame_vm_group_bin_15322 (RW)
0x3b: frame_vm_group_bin_8131 (RW)
0x3c: frame_vm_group_bin_0977 (RW)
0x3d: frame_vm_group_bin_17170 (RW)
0x3e: frame_vm_group_bin_9961 (RW)
0x3f: frame_vm_group_bin_2803 (RW)
0x40: frame_vm_group_bin_18877 (RW)
0x41: frame_vm_group_bin_11749 (RW)
0x42: frame_vm_group_bin_4613 (RW)
0x43: frame_vm_group_bin_20729 (RW)
0x44: frame_vm_group_bin_13530 (RW)
0x45: frame_vm_group_bin_6344 (RW)
0x46: frame_vm_group_bin_22537 (RW)
0x47: frame_vm_group_bin_15355 (RW)
0x48: frame_vm_group_bin_8164 (RW)
0x49: frame_vm_group_bin_1010 (RW)
0x4: frame_vm_group_bin_6189 (RW)
0x4a: frame_vm_group_bin_17201 (RW)
0x4b: frame_vm_group_bin_9994 (RW)
0x4c: frame_vm_group_bin_2836 (RW)
0x4d: frame_vm_group_bin_18910 (RW)
0x4e: frame_vm_group_bin_11772 (RW)
0x4f: frame_vm_group_bin_4641 (RW)
0x50: frame_vm_group_bin_20762 (RW)
0x51: frame_vm_group_bin_13563 (RW)
0x52: frame_vm_group_bin_6376 (RW)
0x53: frame_vm_group_bin_22570 (RW)
0x54: frame_vm_group_bin_15388 (RW)
0x55: frame_vm_group_bin_8197 (RW)
0x56: frame_vm_group_bin_16485 (RW)
0x57: frame_vm_group_bin_17234 (RW)
0x58: frame_vm_group_bin_10027 (RW)
0x59: frame_vm_group_bin_2870 (RW)
0x5: frame_vm_group_bin_22372 (RW)
0x5a: frame_vm_group_bin_18943 (RW)
0x5b: frame_vm_group_bin_11800 (RW)
0x5c: frame_vm_group_bin_4675 (RW)
0x5d: frame_vm_group_bin_20796 (RW)
0x5e: frame_vm_group_bin_13597 (RW)
0x5f: frame_vm_group_bin_6407 (RW)
0x60: frame_vm_group_bin_22604 (RW)
0x61: frame_vm_group_bin_15422 (RW)
0x62: frame_vm_group_bin_8231 (RW)
0x63: frame_vm_group_bin_21118 (RW)
0x64: frame_vm_group_bin_17267 (RW)
0x65: frame_vm_group_bin_10061 (RW)
0x66: frame_vm_group_bin_2904 (RW)
0x67: frame_vm_group_bin_18974 (RW)
0x68: frame_vm_group_bin_11833 (RW)
0x69: frame_vm_group_bin_4706 (RW)
0x6: frame_vm_group_bin_15188 (RW)
0x6a: frame_vm_group_bin_20828 (RW)
0x6b: frame_vm_group_bin_13630 (RW)
0x6c: frame_vm_group_bin_6440 (RW)
0x6d: frame_vm_group_bin_22637 (RW)
0x6e: frame_vm_group_bin_15455 (RW)
0x6f: frame_vm_group_bin_8264 (RW)
0x70: frame_vm_group_bin_1079 (RW)
0x71: frame_vm_group_bin_17300 (RW)
0x72: frame_vm_group_bin_10094 (RW)
0x73: frame_vm_group_bin_2937 (RW)
0x74: frame_vm_group_bin_19007 (RW)
0x75: frame_vm_group_bin_11861 (RW)
0x76: frame_vm_group_bin_4738 (RW)
0x77: frame_vm_group_bin_15771 (RW)
0x78: frame_vm_group_bin_13662 (RW)
0x79: frame_vm_group_bin_6473 (RW)
0x7: frame_vm_group_bin_13168 (RW)
0x7a: frame_vm_group_bin_22671 (RW)
0x7b: frame_vm_group_bin_15489 (RW)
0x7c: frame_vm_group_bin_8297 (RW)
0x7d: frame_vm_group_bin_1109 (RW)
0x7e: frame_vm_group_bin_17334 (RW)
0x7f: frame_vm_group_bin_10128 (RW)
0x80: frame_vm_group_bin_2971 (RW)
0x81: frame_vm_group_bin_19041 (RW)
0x82: frame_vm_group_bin_11889 (RW)
0x83: frame_vm_group_bin_4772 (RW)
0x84: frame_vm_group_bin_20881 (RW)
0x85: frame_vm_group_bin_13696 (RW)
0x86: frame_vm_group_bin_6507 (RW)
0x87: frame_vm_group_bin_22704 (RW)
0x88: frame_vm_group_bin_15521 (RW)
0x89: frame_vm_group_bin_8330 (RW)
0x8: frame_vm_group_bin_0843 (RW)
0x8a: frame_vm_group_bin_1141 (RW)
0x8b: frame_vm_group_bin_17366 (RW)
0x8c: frame_vm_group_bin_10163 (RW)
0x8d: frame_vm_group_bin_3004 (RW)
0x8e: frame_vm_group_bin_19074 (RW)
0x8f: frame_vm_group_bin_11913 (RW)
0x90: frame_vm_group_bin_4805 (RW)
0x91: frame_vm_group_bin_20909 (RW)
0x92: frame_vm_group_bin_13728 (RW)
0x93: frame_vm_group_bin_6540 (RW)
0x94: frame_vm_group_bin_22737 (RW)
0x95: frame_vm_group_bin_15553 (RW)
0x96: frame_vm_group_bin_8363 (RW)
0x97: frame_vm_group_bin_1174 (RW)
0x98: frame_vm_group_bin_17396 (RW)
0x99: frame_vm_group_bin_10196 (RW)
0x9: frame_vm_group_bin_17038 (RW)
0x9a: frame_vm_group_bin_3038 (RW)
0x9b: frame_vm_group_bin_19108 (RW)
0x9c: frame_vm_group_bin_11943 (RW)
0x9d: frame_vm_group_bin_4838 (RW)
0x9e: frame_vm_group_bin_20939 (RW)
0x9f: frame_vm_group_bin_13763 (RW)
0xa0: frame_vm_group_bin_6574 (RW)
0xa1: frame_vm_group_bin_22770 (RW)
0xa2: frame_vm_group_bin_15587 (RW)
0xa3: frame_vm_group_bin_8397 (RW)
0xa4: frame_vm_group_bin_1208 (RW)
0xa5: frame_vm_group_bin_17422 (RW)
0xa6: frame_vm_group_bin_10230 (RW)
0xa7: frame_vm_group_bin_3071 (RW)
0xa8: frame_vm_group_bin_19139 (RW)
0xa9: frame_vm_group_bin_11976 (RW)
0xa: frame_vm_group_bin_9830 (RW)
0xaa: frame_vm_group_bin_4871 (RW)
0xab: frame_vm_group_bin_20964 (RW)
0xac: frame_vm_group_bin_13796 (RW)
0xad: frame_vm_group_bin_6607 (RW)
0xae: frame_vm_group_bin_22803 (RW)
0xaf: frame_vm_group_bin_15620 (RW)
0xb0: frame_vm_group_bin_8430 (RW)
0xb1: frame_vm_group_bin_1241 (RW)
0xb2: frame_vm_group_bin_17447 (RW)
0xb3: frame_vm_group_bin_10263 (RW)
0xb4: frame_vm_group_bin_3104 (RW)
0xb5: frame_vm_group_bin_19172 (RW)
0xb6: frame_vm_group_bin_12008 (RW)
0xb7: frame_vm_group_bin_4904 (RW)
0xb8: frame_vm_group_bin_20997 (RW)
0xb9: frame_vm_group_bin_13827 (RW)
0xb: frame_vm_group_bin_2669 (RW)
0xba: frame_vm_group_bin_6641 (RW)
0xbb: frame_vm_group_bin_22837 (RW)
0xbc: frame_vm_group_bin_15654 (RW)
0xbd: frame_vm_group_bin_8464 (RW)
0xbe: frame_vm_group_bin_1272 (RW)
0xbf: frame_vm_group_bin_17468 (RW)
0xc0: frame_vm_group_bin_10297 (RW)
0xc1: frame_vm_group_bin_3137 (RW)
0xc2: frame_vm_group_bin_19206 (RW)
0xc3: frame_vm_group_bin_12039 (RW)
0xc4: frame_vm_group_bin_4936 (RW)
0xc5: frame_vm_group_bin_21031 (RW)
0xc6: frame_vm_group_bin_13857 (RW)
0xc7: frame_vm_group_bin_6674 (RW)
0xc8: frame_vm_group_bin_22870 (RW)
0xc9: frame_vm_group_bin_15687 (RW)
0xc: frame_vm_group_bin_18742 (RW)
0xca: frame_vm_group_bin_8497 (RW)
0xcb: frame_vm_group_bin_1305 (RW)
0xcc: frame_vm_group_bin_17490 (RW)
0xcd: frame_vm_group_bin_10330 (RW)
0xce: frame_vm_group_bin_3170 (RW)
0xcf: frame_vm_group_bin_19239 (RW)
0xd0: frame_vm_group_bin_12066 (RW)
0xd1: frame_vm_group_bin_4967 (RW)
0xd2: frame_vm_group_bin_21065 (RW)
0xd3: frame_vm_group_bin_13887 (RW)
0xd4: frame_vm_group_bin_6707 (RW)
0xd5: frame_vm_group_bin_22903 (RW)
0xd6: frame_vm_group_bin_15720 (RW)
0xd7: frame_vm_group_bin_8529 (RW)
0xd8: frame_vm_group_bin_1337 (RW)
0xd9: frame_vm_group_bin_17515 (RW)
0xd: frame_vm_group_bin_11651 (RW)
0xda: frame_vm_group_bin_10364 (RW)
0xdb: frame_vm_group_bin_3204 (RW)
0xdc: frame_vm_group_bin_19273 (RW)
0xdd: frame_vm_group_bin_12100 (RW)
0xde: frame_vm_group_bin_5001 (RW)
0xdf: frame_vm_group_bin_21099 (RW)
0xe0: frame_vm_group_bin_13921 (RW)
0xe1: frame_vm_group_bin_6740 (RW)
0xe2: frame_vm_group_bin_22937 (RW)
0xe3: frame_vm_group_bin_15754 (RW)
0xe4: frame_vm_group_bin_8561 (RW)
0xe5: frame_vm_group_bin_1372 (RW)
0xe6: frame_vm_group_bin_17542 (RW)
0xe7: frame_vm_group_bin_18260 (RW)
0xe8: frame_vm_group_bin_3236 (RW)
0xe9: frame_vm_group_bin_19306 (RW)
0xe: frame_vm_group_bin_4500 (RW)
0xea: frame_vm_group_bin_12132 (RW)
0xeb: frame_vm_group_bin_5034 (RW)
0xec: frame_vm_group_bin_21132 (RW)
0xed: frame_vm_group_bin_13954 (RW)
0xee: frame_vm_group_bin_6772 (RW)
0xef: frame_vm_group_bin_22969 (RW)
0xf0: frame_vm_group_bin_15787 (RW)
0xf1: frame_vm_group_bin_8594 (RW)
0xf2: frame_vm_group_bin_1405 (RW)
0xf3: frame_vm_group_bin_17563 (RW)
0xf4: frame_vm_group_bin_10419 (RW)
0xf5: frame_vm_group_bin_3269 (RW)
0xf6: frame_vm_group_bin_19339 (RW)
0xf7: frame_vm_group_bin_18614 (RW)
0xf8: frame_vm_group_bin_5067 (RW)
0xf9: frame_vm_group_bin_21164 (RW)
0xf: frame_vm_group_bin_20596 (RW)
0xfa: frame_vm_group_bin_13988 (RW)
0xfb: frame_vm_group_bin_6806 (RW)
0xfc: frame_vm_group_bin_23002 (RW)
0xfd: frame_vm_group_bin_10076 (RW)
0xfe: frame_vm_group_bin_8627 (RW)
0xff: frame_vm_group_bin_1439 (RW)
}
pt_vm_group_bin_0060 {
0x0: frame_vm_group_bin_1747 (RW)
0x100: frame_vm_group_bin_7743 (RW)
0x101: frame_vm_group_bin_0580 (RW)
0x102: frame_vm_group_bin_16774 (RW)
0x103: frame_vm_group_bin_9565 (RW)
0x104: frame_vm_group_bin_2405 (RW)
0x105: frame_vm_group_bin_18497 (RW)
0x106: frame_vm_group_bin_11416 (RW)
0x107: frame_vm_group_bin_4232 (RW)
0x108: frame_vm_group_bin_20330 (RW)
0x109: frame_vm_group_bin_13133 (RW)
0x10: frame_vm_group_bin_3602 (RW)
0x10a: frame_vm_group_bin_5980 (RW)
0x10b: frame_vm_group_bin_22141 (RW)
0x10c: frame_vm_group_bin_14992 (RW)
0x10d: frame_vm_group_bin_7776 (RW)
0x10e: frame_vm_group_bin_0612 (RW)
0x10f: frame_vm_group_bin_16807 (RW)
0x110: frame_vm_group_bin_9598 (RW)
0x111: frame_vm_group_bin_2437 (RW)
0x112: frame_vm_group_bin_18523 (RW)
0x113: frame_vm_group_bin_11449 (RW)
0x114: frame_vm_group_bin_4265 (RW)
0x115: frame_vm_group_bin_20363 (RW)
0x116: frame_vm_group_bin_13166 (RW)
0x117: frame_vm_group_bin_6011 (RW)
0x118: frame_vm_group_bin_22174 (RW)
0x119: frame_vm_group_bin_15025 (RW)
0x11: frame_vm_group_bin_19702 (RW)
0x11a: frame_vm_group_bin_7810 (RW)
0x11b: frame_vm_group_bin_0645 (RW)
0x11c: frame_vm_group_bin_16841 (RW)
0x11d: frame_vm_group_bin_9632 (RW)
0x11e: frame_vm_group_bin_2470 (RW)
0x11f: frame_vm_group_bin_18551 (RW)
0x120: frame_vm_group_bin_11483 (RW)
0x121: frame_vm_group_bin_4299 (RW)
0x122: frame_vm_group_bin_20397 (RW)
0x123: frame_vm_group_bin_13200 (RW)
0x124: frame_vm_group_bin_6042 (RW)
0x125: frame_vm_group_bin_22208 (RW)
0x126: frame_vm_group_bin_9533 (RW)
0x127: frame_vm_group_bin_7842 (RW)
0x128: frame_vm_group_bin_0678 (RW)
0x129: frame_vm_group_bin_16873 (RW)
0x12: frame_vm_group_bin_12530 (RW)
0x12a: frame_vm_group_bin_9665 (RW)
0x12b: frame_vm_group_bin_2503 (RW)
0x12c: frame_vm_group_bin_18580 (RW)
0x12d: frame_vm_group_bin_11516 (RW)
0x12e: frame_vm_group_bin_4332 (RW)
0x12f: frame_vm_group_bin_20430 (RW)
0x130: frame_vm_group_bin_13233 (RW)
0x131: frame_vm_group_bin_6065 (RW)
0x132: frame_vm_group_bin_22241 (RW)
0x133: frame_vm_group_bin_15075 (RW)
0x134: frame_vm_group_bin_7875 (RW)
0x135: frame_vm_group_bin_0711 (RW)
0x136: frame_vm_group_bin_16905 (RW)
0x137: frame_vm_group_bin_9697 (RW)
0x138: frame_vm_group_bin_2536 (RW)
0x139: frame_vm_group_bin_18613 (RW)
0x13: frame_vm_group_bin_5440 (RW)
0x13a: frame_vm_group_bin_11550 (RW)
0x13b: frame_vm_group_bin_4368 (RW)
0x13c: frame_vm_group_bin_20464 (RW)
0x13d: frame_vm_group_bin_13267 (RW)
0x13e: frame_vm_group_bin_6094 (RW)
0x13f: frame_vm_group_bin_22274 (RW)
0x140: frame_vm_group_bin_15103 (RW)
0x141: frame_vm_group_bin_7909 (RW)
0x142: frame_vm_group_bin_0745 (RW)
0x143: frame_vm_group_bin_16939 (RW)
0x144: frame_vm_group_bin_9731 (RW)
0x145: frame_vm_group_bin_2570 (RW)
0x146: frame_vm_group_bin_18646 (RW)
0x147: frame_vm_group_bin_11578 (RW)
0x148: frame_vm_group_bin_4401 (RW)
0x149: frame_vm_group_bin_20497 (RW)
0x14: frame_vm_group_bin_21535 (RW)
0x14a: frame_vm_group_bin_13300 (RW)
0x14b: frame_vm_group_bin_6125 (RW)
0x14c: frame_vm_group_bin_22307 (RW)
0x14d: frame_vm_group_bin_15129 (RW)
0x14e: frame_vm_group_bin_7943 (RW)
0x14f: frame_vm_group_bin_0778 (RW)
0x150: frame_vm_group_bin_16972 (RW)
0x151: frame_vm_group_bin_9764 (RW)
0x152: frame_vm_group_bin_2603 (RW)
0x153: frame_vm_group_bin_18679 (RW)
0x154: frame_vm_group_bin_11602 (RW)
0x155: frame_vm_group_bin_4434 (RW)
0x156: frame_vm_group_bin_20530 (RW)
0x157: frame_vm_group_bin_13332 (RW)
0x158: frame_vm_group_bin_6157 (RW)
0x159: frame_vm_group_bin_22339 (RW)
0x15: frame_vm_group_bin_14359 (RW)
0x15a: frame_vm_group_bin_15156 (RW)
0x15b: frame_vm_group_bin_7977 (RW)
0x15c: frame_vm_group_bin_0811 (RW)
0x15d: frame_vm_group_bin_17006 (RW)
0x15e: frame_vm_group_bin_9798 (RW)
0x15f: frame_vm_group_bin_2637 (RW)
0x160: frame_vm_group_bin_18712 (RW)
0x161: frame_vm_group_bin_11630 (RW)
0x162: frame_vm_group_bin_4468 (RW)
0x163: frame_vm_group_bin_20564 (RW)
0x164: frame_vm_group_bin_13366 (RW)
0x165: frame_vm_group_bin_6190 (RW)
0x166: frame_vm_group_bin_22373 (RW)
0x167: frame_vm_group_bin_15189 (RW)
0x168: frame_vm_group_bin_8007 (RW)
0x169: frame_vm_group_bin_0844 (RW)
0x16: frame_vm_group_bin_7144 (RW)
0x16a: frame_vm_group_bin_17039 (RW)
0x16b: frame_vm_group_bin_9831 (RW)
0x16c: frame_vm_group_bin_2670 (RW)
0x16d: frame_vm_group_bin_18743 (RW)
0x16e: frame_vm_group_bin_11652 (RW)
0x16f: frame_vm_group_bin_4501 (RW)
0x170: frame_vm_group_bin_20597 (RW)
0x171: frame_vm_group_bin_13397 (RW)
0x172: frame_vm_group_bin_6217 (RW)
0x173: frame_vm_group_bin_22406 (RW)
0x174: frame_vm_group_bin_15222 (RW)
0x175: frame_vm_group_bin_8035 (RW)
0x176: frame_vm_group_bin_0877 (RW)
0x177: frame_vm_group_bin_17072 (RW)
0x178: frame_vm_group_bin_9864 (RW)
0x179: frame_vm_group_bin_2703 (RW)
0x17: frame_vm_group_bin_0062 (RW)
0x17a: frame_vm_group_bin_18777 (RW)
0x17b: frame_vm_group_bin_11673 (RW)
0x17c: frame_vm_group_bin_4535 (RW)
0x17d: frame_vm_group_bin_20631 (RW)
0x17e: frame_vm_group_bin_13431 (RW)
0x17f: frame_vm_group_bin_6247 (RW)
0x180: frame_vm_group_bin_22439 (RW)
0x181: frame_vm_group_bin_15257 (RW)
0x182: frame_vm_group_bin_8067 (RW)
0x183: frame_vm_group_bin_0911 (RW)
0x184: frame_vm_group_bin_17106 (RW)
0x185: frame_vm_group_bin_9897 (RW)
0x186: frame_vm_group_bin_2737 (RW)
0x187: frame_vm_group_bin_18810 (RW)
0x188: frame_vm_group_bin_11700 (RW)
0x189: frame_vm_group_bin_7385 (RW)
0x18: frame_vm_group_bin_16193 (RW)
0x18a: frame_vm_group_bin_20663 (RW)
0x18b: frame_vm_group_bin_13464 (RW)
0x18c: frame_vm_group_bin_6279 (RW)
0x18d: frame_vm_group_bin_22472 (RW)
0x18e: frame_vm_group_bin_15289 (RW)
0x18f: frame_vm_group_bin_8099 (RW)
0x190: frame_vm_group_bin_0944 (RW)
0x191: frame_vm_group_bin_17139 (RW)
0x192: frame_vm_group_bin_9930 (RW)
0x193: frame_vm_group_bin_2770 (RW)
0x194: frame_vm_group_bin_18844 (RW)
0x195: frame_vm_group_bin_11727 (RW)
0x196: frame_vm_group_bin_4589 (RW)
0x197: frame_vm_group_bin_20696 (RW)
0x198: frame_vm_group_bin_13497 (RW)
0x199: frame_vm_group_bin_6312 (RW)
0x19: frame_vm_group_bin_9000 (RW)
0x19a: frame_vm_group_bin_22506 (RW)
0x19b: frame_vm_group_bin_15323 (RW)
0x19c: frame_vm_group_bin_8132 (RW)
0x19d: frame_vm_group_bin_0978 (RW)
0x19e: frame_vm_group_bin_17171 (RW)
0x19f: frame_vm_group_bin_9962 (RW)
0x1: frame_vm_group_bin_17856 (RW)
0x1a0: frame_vm_group_bin_2804 (RW)
0x1a1: frame_vm_group_bin_18878 (RW)
0x1a2: frame_vm_group_bin_11750 (RW)
0x1a3: frame_vm_group_bin_4614 (RW)
0x1a4: frame_vm_group_bin_20730 (RW)
0x1a5: frame_vm_group_bin_13531 (RW)
0x1a6: frame_vm_group_bin_6345 (RW)
0x1a7: frame_vm_group_bin_22538 (RW)
0x1a8: frame_vm_group_bin_15356 (RW)
0x1a9: frame_vm_group_bin_8165 (RW)
0x1a: frame_vm_group_bin_1813 (RW)
0x1aa: frame_vm_group_bin_6687 (RW)
0x1ab: frame_vm_group_bin_17202 (RW)
0x1ac: frame_vm_group_bin_9995 (RW)
0x1ad: frame_vm_group_bin_2837 (RW)
0x1ae: frame_vm_group_bin_18911 (RW)
0x1af: frame_vm_group_bin_11773 (RW)
0x1b0: frame_vm_group_bin_4642 (RW)
0x1b1: frame_vm_group_bin_20763 (RW)
0x1b2: frame_vm_group_bin_13564 (RW)
0x1b3: frame_vm_group_bin_6377 (RW)
0x1b4: frame_vm_group_bin_22571 (RW)
0x1b5: frame_vm_group_bin_15389 (RW)
0x1b6: frame_vm_group_bin_8198 (RW)
0x1b7: frame_vm_group_bin_1034 (RW)
0x1b8: frame_vm_group_bin_9956 (RW)
0x1b9: frame_vm_group_bin_10028 (RW)
0x1b: frame_vm_group_bin_17915 (RW)
0x1ba: frame_vm_group_bin_2872 (RW)
0x1bb: frame_vm_group_bin_18944 (RW)
0x1bc: frame_vm_group_bin_11801 (RW)
0x1bd: frame_vm_group_bin_2797 (RW)
0x1be: frame_vm_group_bin_20797 (RW)
0x1bf: frame_vm_group_bin_13598 (RW)
0x1c0: frame_vm_group_bin_6408 (RW)
0x1c1: frame_vm_group_bin_22605 (RW)
0x1c2: frame_vm_group_bin_15423 (RW)
0x1c3: frame_vm_group_bin_8232 (RW)
0x1c4: frame_vm_group_bin_1056 (RW)
0x1c5: frame_vm_group_bin_17268 (RW)
0x1c6: frame_vm_group_bin_10062 (RW)
0x1c7: frame_vm_group_bin_2905 (RW)
0x1c8: frame_vm_group_bin_18975 (RW)
0x1c9: frame_vm_group_bin_11834 (RW)
0x1c: frame_vm_group_bin_10821 (RW)
0x1ca: frame_vm_group_bin_4707 (RW)
0x1cb: frame_vm_group_bin_20829 (RW)
0x1cc: frame_vm_group_bin_13631 (RW)
0x1cd: frame_vm_group_bin_6441 (RW)
0x1ce: frame_vm_group_bin_22638 (RW)
0x1cf: frame_vm_group_bin_15456 (RW)
0x1d0: frame_vm_group_bin_8265 (RW)
0x1d1: frame_vm_group_bin_1080 (RW)
0x1d2: frame_vm_group_bin_17301 (RW)
0x1d3: frame_vm_group_bin_10095 (RW)
0x1d4: frame_vm_group_bin_2938 (RW)
0x1d5: frame_vm_group_bin_19008 (RW)
0x1d6: frame_vm_group_bin_11862 (RW)
0x1d7: frame_vm_group_bin_4739 (RW)
0x1d8: frame_vm_group_bin_20857 (RW)
0x1d9: frame_vm_group_bin_13663 (RW)
0x1d: frame_vm_group_bin_3636 (RW)
0x1da: frame_vm_group_bin_6475 (RW)
0x1db: frame_vm_group_bin_22672 (RW)
0x1dc: frame_vm_group_bin_15490 (RW)
0x1dd: frame_vm_group_bin_8298 (RW)
0x1de: frame_vm_group_bin_1110 (RW)
0x1df: frame_vm_group_bin_17335 (RW)
0x1e0: frame_vm_group_bin_10129 (RW)
0x1e1: frame_vm_group_bin_2972 (RW)
0x1e2: frame_vm_group_bin_19042 (RW)
0x1e3: frame_vm_group_bin_11890 (RW)
0x1e4: frame_vm_group_bin_4773 (RW)
0x1e5: frame_vm_group_bin_20882 (RW)
0x1e6: frame_vm_group_bin_13697 (RW)
0x1e7: frame_vm_group_bin_6508 (RW)
0x1e8: frame_vm_group_bin_22705 (RW)
0x1e9: frame_vm_group_bin_15522 (RW)
0x1e: frame_vm_group_bin_19736 (RW)
0x1ea: frame_vm_group_bin_8331 (RW)
0x1eb: frame_vm_group_bin_1142 (RW)
0x1ec: frame_vm_group_bin_17367 (RW)
0x1ed: frame_vm_group_bin_10164 (RW)
0x1ee: frame_vm_group_bin_3005 (RW)
0x1ef: frame_vm_group_bin_19075 (RW)
0x1f0: frame_vm_group_bin_11914 (RW)
0x1f1: frame_vm_group_bin_4806 (RW)
0x1f2: frame_vm_group_bin_20910 (RW)
0x1f3: frame_vm_group_bin_13729 (RW)
0x1f4: frame_vm_group_bin_6541 (RW)
0x1f5: frame_vm_group_bin_22738 (RW)
0x1f6: frame_vm_group_bin_15554 (RW)
0x1f7: frame_vm_group_bin_8364 (RW)
0x1f8: frame_vm_group_bin_1175 (RW)
0x1f9: frame_vm_group_bin_17397 (RW)
0x1f: frame_vm_group_bin_12564 (RW)
0x1fa: frame_vm_group_bin_10198 (RW)
0x1fb: frame_vm_group_bin_3039 (RW)
0x1fc: frame_vm_group_bin_5723 (RW)
0x1fd: frame_vm_group_bin_11944 (RW)
0x1fe: frame_vm_group_bin_4839 (RW)
0x1ff: frame_vm_group_bin_20940 (RW)
0x20: frame_vm_group_bin_5472 (RW)
0x21: frame_vm_group_bin_21569 (RW)
0x22: frame_vm_group_bin_14393 (RW)
0x23: frame_vm_group_bin_7180 (RW)
0x24: frame_vm_group_bin_0089 (RW)
0x25: frame_vm_group_bin_5188 (RW)
0x26: frame_vm_group_bin_9034 (RW)
0x27: frame_vm_group_bin_1846 (RW)
0x28: frame_vm_group_bin_17947 (RW)
0x29: frame_vm_group_bin_10854 (RW)
0x2: frame_vm_group_bin_10755 (RW)
0x2a: frame_vm_group_bin_3669 (RW)
0x2b: frame_vm_group_bin_19769 (RW)
0x2c: frame_vm_group_bin_12597 (RW)
0x2d: frame_vm_group_bin_5505 (RW)
0x2e: frame_vm_group_bin_21602 (RW)
0x2f: frame_vm_group_bin_14426 (RW)
0x30: frame_vm_group_bin_7213 (RW)
0x31: frame_vm_group_bin_0114 (RW)
0x32: frame_vm_group_bin_16247 (RW)
0x33: frame_vm_group_bin_9067 (RW)
0x34: frame_vm_group_bin_1879 (RW)
0x35: frame_vm_group_bin_17977 (RW)
0x36: frame_vm_group_bin_10886 (RW)
0x37: frame_vm_group_bin_3702 (RW)
0x38: frame_vm_group_bin_19802 (RW)
0x39: frame_vm_group_bin_12630 (RW)
0x3: frame_vm_group_bin_3568 (RW)
0x3a: frame_vm_group_bin_5538 (RW)
0x3b: frame_vm_group_bin_21636 (RW)
0x3c: frame_vm_group_bin_14460 (RW)
0x3d: frame_vm_group_bin_7247 (RW)
0x3e: frame_vm_group_bin_0137 (RW)
0x3f: frame_vm_group_bin_16278 (RW)
0x40: frame_vm_group_bin_9101 (RW)
0x41: frame_vm_group_bin_1913 (RW)
0x42: frame_vm_group_bin_18011 (RW)
0x43: frame_vm_group_bin_10921 (RW)
0x44: frame_vm_group_bin_3736 (RW)
0x45: frame_vm_group_bin_19836 (RW)
0x46: frame_vm_group_bin_4486 (RW)
0x47: frame_vm_group_bin_5571 (RW)
0x48: frame_vm_group_bin_21669 (RW)
0x49: frame_vm_group_bin_14493 (RW)
0x4: frame_vm_group_bin_19672 (RW)
0x4a: frame_vm_group_bin_7280 (RW)
0x4b: frame_vm_group_bin_0158 (RW)
0x4c: frame_vm_group_bin_16309 (RW)
0x4d: frame_vm_group_bin_9134 (RW)
0x4e: frame_vm_group_bin_1946 (RW)
0x4f: frame_vm_group_bin_18044 (RW)
0x50: frame_vm_group_bin_10954 (RW)
0x51: frame_vm_group_bin_3769 (RW)
0x52: frame_vm_group_bin_19869 (RW)
0x53: frame_vm_group_bin_12683 (RW)
0x54: frame_vm_group_bin_5603 (RW)
0x55: frame_vm_group_bin_21701 (RW)
0x56: frame_vm_group_bin_14527 (RW)
0x57: frame_vm_group_bin_7312 (RW)
0x58: frame_vm_group_bin_0187 (RW)
0x59: frame_vm_group_bin_16341 (RW)
0x5: frame_vm_group_bin_12497 (RW)
0x5a: frame_vm_group_bin_9166 (RW)
0x5b: frame_vm_group_bin_1979 (RW)
0x5c: frame_vm_group_bin_19480 (RW)
0x5d: frame_vm_group_bin_10987 (RW)
0x5e: frame_vm_group_bin_3802 (RW)
0x5f: frame_vm_group_bin_19901 (RW)
0x60: frame_vm_group_bin_12711 (RW)
0x61: frame_vm_group_bin_5635 (RW)
0x62: frame_vm_group_bin_21735 (RW)
0x63: frame_vm_group_bin_14561 (RW)
0x64: frame_vm_group_bin_7346 (RW)
0x65: frame_vm_group_bin_0219 (RW)
0x66: frame_vm_group_bin_16375 (RW)
0x67: frame_vm_group_bin_3752 (RW)
0x68: frame_vm_group_bin_2012 (RW)
0x69: frame_vm_group_bin_18108 (RW)
0x6: frame_vm_group_bin_5407 (RW)
0x6a: frame_vm_group_bin_11020 (RW)
0x6b: frame_vm_group_bin_3835 (RW)
0x6c: frame_vm_group_bin_19933 (RW)
0x6d: frame_vm_group_bin_12735 (RW)
0x6e: frame_vm_group_bin_5668 (RW)
0x6f: frame_vm_group_bin_21768 (RW)
0x70: frame_vm_group_bin_14594 (RW)
0x71: frame_vm_group_bin_7379 (RW)
0x72: frame_vm_group_bin_0244 (RW)
0x73: frame_vm_group_bin_16408 (RW)
0x74: frame_vm_group_bin_9222 (RW)
0x75: frame_vm_group_bin_2045 (RW)
0x76: frame_vm_group_bin_18141 (RW)
0x77: frame_vm_group_bin_11053 (RW)
0x78: frame_vm_group_bin_3868 (RW)
0x79: frame_vm_group_bin_19966 (RW)
0x7: frame_vm_group_bin_21502 (RW)
0x7a: frame_vm_group_bin_12766 (RW)
0x7b: frame_vm_group_bin_5702 (RW)
0x7c: frame_vm_group_bin_21802 (RW)
0x7d: frame_vm_group_bin_14627 (RW)
0x7e: frame_vm_group_bin_7413 (RW)
0x7f: frame_vm_group_bin_0267 (RW)
0x80: frame_vm_group_bin_16442 (RW)
0x81: frame_vm_group_bin_9248 (RW)
0x82: frame_vm_group_bin_2079 (RW)
0x83: frame_vm_group_bin_18175 (RW)
0x84: frame_vm_group_bin_11087 (RW)
0x85: frame_vm_group_bin_3902 (RW)
0x86: frame_vm_group_bin_19998 (RW)
0x87: frame_vm_group_bin_12799 (RW)
0x88: frame_vm_group_bin_3060 (RW)
0x89: frame_vm_group_bin_21835 (RW)
0x8: frame_vm_group_bin_14326 (RW)
0x8a: frame_vm_group_bin_14660 (RW)
0x8b: frame_vm_group_bin_7446 (RW)
0x8c: frame_vm_group_bin_0294 (RW)
0x8d: frame_vm_group_bin_16475 (RW)
0x8e: frame_vm_group_bin_9270 (RW)
0x8f: frame_vm_group_bin_2112 (RW)
0x90: frame_vm_group_bin_18207 (RW)
0x91: frame_vm_group_bin_11120 (RW)
0x92: frame_vm_group_bin_3935 (RW)
0x93: frame_vm_group_bin_20031 (RW)
0x94: frame_vm_group_bin_12831 (RW)
0x95: frame_vm_group_bin_5759 (RW)
0x96: frame_vm_group_bin_21868 (RW)
0x97: frame_vm_group_bin_14693 (RW)
0x98: frame_vm_group_bin_7479 (RW)
0x99: frame_vm_group_bin_0326 (RW)
0x9: frame_vm_group_bin_7112 (RW)
0x9a: frame_vm_group_bin_16509 (RW)
0x9b: frame_vm_group_bin_22410 (RW)
0x9c: frame_vm_group_bin_2147 (RW)
0x9d: frame_vm_group_bin_18241 (RW)
0x9e: frame_vm_group_bin_11153 (RW)
0x9f: frame_vm_group_bin_3968 (RW)
0xa0: frame_vm_group_bin_20065 (RW)
0xa1: frame_vm_group_bin_12865 (RW)
0xa2: frame_vm_group_bin_5784 (RW)
0xa3: frame_vm_group_bin_21902 (RW)
0xa4: frame_vm_group_bin_14727 (RW)
0xa5: frame_vm_group_bin_7512 (RW)
0xa6: frame_vm_group_bin_0358 (RW)
0xa7: frame_vm_group_bin_16542 (RW)
0xa8: frame_vm_group_bin_9330 (RW)
0xa9: frame_vm_group_bin_2180 (RW)
0xa: frame_vm_group_bin_0037 (RW)
0xaa: frame_vm_group_bin_18274 (RW)
0xab: frame_vm_group_bin_11186 (RW)
0xac: frame_vm_group_bin_4001 (RW)
0xad: frame_vm_group_bin_20098 (RW)
0xae: frame_vm_group_bin_12898 (RW)
0xaf: frame_vm_group_bin_5806 (RW)
0xb0: frame_vm_group_bin_21934 (RW)
0xb1: frame_vm_group_bin_14759 (RW)
0xb2: frame_vm_group_bin_7544 (RW)
0xb3: frame_vm_group_bin_0389 (RW)
0xb4: frame_vm_group_bin_16574 (RW)
0xb5: frame_vm_group_bin_9363 (RW)
0xb6: frame_vm_group_bin_2209 (RW)
0xb7: frame_vm_group_bin_18307 (RW)
0xb8: frame_vm_group_bin_11219 (RW)
0xb9: frame_vm_group_bin_4034 (RW)
0xb: frame_vm_group_bin_16160 (RW)
0xba: frame_vm_group_bin_20131 (RW)
0xbb: frame_vm_group_bin_12931 (RW)
0xbc: frame_vm_group_bin_5829 (RW)
0xbd: frame_vm_group_bin_21968 (RW)
0xbe: frame_vm_group_bin_14792 (RW)
0xbf: frame_vm_group_bin_7577 (RW)
0xc0: frame_vm_group_bin_0418 (RW)
0xc1: frame_vm_group_bin_16607 (RW)
0xc2: frame_vm_group_bin_9398 (RW)
0xc3: frame_vm_group_bin_2239 (RW)
0xc4: frame_vm_group_bin_18341 (RW)
0xc5: frame_vm_group_bin_11253 (RW)
0xc6: frame_vm_group_bin_4068 (RW)
0xc7: frame_vm_group_bin_20163 (RW)
0xc8: frame_vm_group_bin_12964 (RW)
0xc9: frame_vm_group_bin_5853 (RW)
0xc: frame_vm_group_bin_8967 (RW)
0xca: frame_vm_group_bin_22001 (RW)
0xcb: frame_vm_group_bin_14825 (RW)
0xcc: frame_vm_group_bin_7610 (RW)
0xcd: frame_vm_group_bin_0450 (RW)
0xce: frame_vm_group_bin_16640 (RW)
0xcf: frame_vm_group_bin_9431 (RW)
0xd0: frame_vm_group_bin_2271 (RW)
0xd1: frame_vm_group_bin_18374 (RW)
0xd2: frame_vm_group_bin_11286 (RW)
0xd3: frame_vm_group_bin_4101 (RW)
0xd4: frame_vm_group_bin_20195 (RW)
0xd5: frame_vm_group_bin_12997 (RW)
0xd6: frame_vm_group_bin_5879 (RW)
0xd7: frame_vm_group_bin_6242 (RW)
0xd8: frame_vm_group_bin_14858 (RW)
0xd9: frame_vm_group_bin_7643 (RW)
0xd: frame_vm_group_bin_1779 (RW)
0xda: frame_vm_group_bin_1977 (RW)
0xdb: frame_vm_group_bin_16674 (RW)
0xdc: frame_vm_group_bin_9465 (RW)
0xdd: frame_vm_group_bin_2305 (RW)
0xde: frame_vm_group_bin_18406 (RW)
0xdf: frame_vm_group_bin_11320 (RW)
0xe0: frame_vm_group_bin_4134 (RW)
0xe1: frame_vm_group_bin_20229 (RW)
0xe2: frame_vm_group_bin_13033 (RW)
0xe3: frame_vm_group_bin_5906 (RW)
0xe4: frame_vm_group_bin_22050 (RW)
0xe5: frame_vm_group_bin_14892 (RW)
0xe6: frame_vm_group_bin_7677 (RW)
0xe7: frame_vm_group_bin_0516 (RW)
0xe8: frame_vm_group_bin_16706 (RW)
0xe9: frame_vm_group_bin_9498 (RW)
0xe: frame_vm_group_bin_17883 (RW)
0xea: frame_vm_group_bin_2338 (RW)
0xeb: frame_vm_group_bin_18439 (RW)
0xec: frame_vm_group_bin_11351 (RW)
0xed: frame_vm_group_bin_4166 (RW)
0xee: frame_vm_group_bin_20262 (RW)
0xef: frame_vm_group_bin_13066 (RW)
0xf0: frame_vm_group_bin_5931 (RW)
0xf1: frame_vm_group_bin_22076 (RW)
0xf2: frame_vm_group_bin_14925 (RW)
0xf3: frame_vm_group_bin_7710 (RW)
0xf4: frame_vm_group_bin_0548 (RW)
0xf5: frame_vm_group_bin_16740 (RW)
0xf6: frame_vm_group_bin_9531 (RW)
0xf7: frame_vm_group_bin_2371 (RW)
0xf8: frame_vm_group_bin_18470 (RW)
0xf9: frame_vm_group_bin_11383 (RW)
0xf: frame_vm_group_bin_10787 (RW)
0xfa: frame_vm_group_bin_4199 (RW)
0xfb: frame_vm_group_bin_20295 (RW)
0xfc: frame_vm_group_bin_13100 (RW)
0xfd: frame_vm_group_bin_5953 (RW)
0xfe: frame_vm_group_bin_22108 (RW)
0xff: frame_vm_group_bin_14959 (RW)
}
pt_vm_group_bin_0063 {
0x0: frame_vm_group_bin_11924 (RW)
0x100: frame_vm_group_bin_17917 (RW)
0x101: frame_vm_group_bin_10823 (RW)
0x102: frame_vm_group_bin_3638 (RW)
0x103: frame_vm_group_bin_19738 (RW)
0x104: frame_vm_group_bin_12566 (RW)
0x105: frame_vm_group_bin_5474 (RW)
0x106: frame_vm_group_bin_21571 (RW)
0x107: frame_vm_group_bin_14395 (RW)
0x108: frame_vm_group_bin_7182 (RW)
0x109: frame_vm_group_bin_4554 (RW)
0x10: frame_vm_group_bin_13774 (RW)
0x10a: frame_vm_group_bin_16223 (RW)
0x10b: frame_vm_group_bin_9036 (RW)
0x10c: frame_vm_group_bin_1848 (RW)
0x10d: frame_vm_group_bin_17949 (RW)
0x10e: frame_vm_group_bin_10856 (RW)
0x10f: frame_vm_group_bin_3671 (RW)
0x110: frame_vm_group_bin_19771 (RW)
0x111: frame_vm_group_bin_12599 (RW)
0x112: frame_vm_group_bin_5507 (RW)
0x113: frame_vm_group_bin_21604 (RW)
0x114: frame_vm_group_bin_14428 (RW)
0x115: frame_vm_group_bin_7215 (RW)
0x116: frame_vm_group_bin_9187 (RW)
0x117: frame_vm_group_bin_16249 (RW)
0x118: frame_vm_group_bin_9069 (RW)
0x119: frame_vm_group_bin_1881 (RW)
0x11: frame_vm_group_bin_6585 (RW)
0x11a: frame_vm_group_bin_17980 (RW)
0x11b: frame_vm_group_bin_10890 (RW)
0x11c: frame_vm_group_bin_3705 (RW)
0x11d: frame_vm_group_bin_19805 (RW)
0x11e: frame_vm_group_bin_12633 (RW)
0x11f: frame_vm_group_bin_5540 (RW)
0x120: frame_vm_group_bin_21638 (RW)
0x121: frame_vm_group_bin_14462 (RW)
0x122: frame_vm_group_bin_7249 (RW)
0x123: frame_vm_group_bin_13828 (RW)
0x124: frame_vm_group_bin_16280 (RW)
0x125: frame_vm_group_bin_9103 (RW)
0x126: frame_vm_group_bin_1915 (RW)
0x127: frame_vm_group_bin_18013 (RW)
0x128: frame_vm_group_bin_10923 (RW)
0x129: frame_vm_group_bin_3738 (RW)
0x12: frame_vm_group_bin_22781 (RW)
0x12a: frame_vm_group_bin_19838 (RW)
0x12b: frame_vm_group_bin_12662 (RW)
0x12c: frame_vm_group_bin_5573 (RW)
0x12d: frame_vm_group_bin_21671 (RW)
0x12e: frame_vm_group_bin_14495 (RW)
0x12f: frame_vm_group_bin_7282 (RW)
0x130: frame_vm_group_bin_18472 (RW)
0x131: frame_vm_group_bin_16311 (RW)
0x132: frame_vm_group_bin_9136 (RW)
0x133: frame_vm_group_bin_1948 (RW)
0x134: frame_vm_group_bin_18046 (RW)
0x135: frame_vm_group_bin_10956 (RW)
0x136: frame_vm_group_bin_3771 (RW)
0x137: frame_vm_group_bin_19871 (RW)
0x138: frame_vm_group_bin_12685 (RW)
0x139: frame_vm_group_bin_5605 (RW)
0x13: frame_vm_group_bin_15598 (RW)
0x13a: frame_vm_group_bin_21704 (RW)
0x13b: frame_vm_group_bin_14530 (RW)
0x13c: frame_vm_group_bin_7315 (RW)
0x13d: frame_vm_group_bin_0190 (RW)
0x13e: frame_vm_group_bin_16344 (RW)
0x13f: frame_vm_group_bin_9168 (RW)
0x140: frame_vm_group_bin_1981 (RW)
0x141: frame_vm_group_bin_18078 (RW)
0x142: frame_vm_group_bin_10989 (RW)
0x143: frame_vm_group_bin_3804 (RW)
0x144: frame_vm_group_bin_19903 (RW)
0x145: frame_vm_group_bin_12713 (RW)
0x146: frame_vm_group_bin_5637 (RW)
0x147: frame_vm_group_bin_21737 (RW)
0x148: frame_vm_group_bin_14563 (RW)
0x149: frame_vm_group_bin_7348 (RW)
0x14: frame_vm_group_bin_8408 (RW)
0x14a: frame_vm_group_bin_4574 (RW)
0x14b: frame_vm_group_bin_16377 (RW)
0x14c: frame_vm_group_bin_9199 (RW)
0x14d: frame_vm_group_bin_2014 (RW)
0x14e: frame_vm_group_bin_18110 (RW)
0x14f: frame_vm_group_bin_11022 (RW)
0x150: frame_vm_group_bin_3837 (RW)
0x151: frame_vm_group_bin_19935 (RW)
0x152: frame_vm_group_bin_12737 (RW)
0x153: frame_vm_group_bin_5670 (RW)
0x154: frame_vm_group_bin_21770 (RW)
0x155: frame_vm_group_bin_14596 (RW)
0x156: frame_vm_group_bin_7381 (RW)
0x157: frame_vm_group_bin_9207 (RW)
0x158: frame_vm_group_bin_16410 (RW)
0x159: frame_vm_group_bin_9224 (RW)
0x15: frame_vm_group_bin_1219 (RW)
0x15a: frame_vm_group_bin_2048 (RW)
0x15b: frame_vm_group_bin_18144 (RW)
0x15c: frame_vm_group_bin_11056 (RW)
0x15d: frame_vm_group_bin_3871 (RW)
0x15e: frame_vm_group_bin_19969 (RW)
0x15f: frame_vm_group_bin_12768 (RW)
0x160: frame_vm_group_bin_5704 (RW)
0x161: frame_vm_group_bin_21804 (RW)
0x162: frame_vm_group_bin_14629 (RW)
0x163: frame_vm_group_bin_7415 (RW)
0x164: frame_vm_group_bin_13848 (RW)
0x165: frame_vm_group_bin_16444 (RW)
0x166: frame_vm_group_bin_9250 (RW)
0x167: frame_vm_group_bin_2081 (RW)
0x168: frame_vm_group_bin_18177 (RW)
0x169: frame_vm_group_bin_11089 (RW)
0x16: frame_vm_group_bin_17430 (RW)
0x16a: frame_vm_group_bin_3904 (RW)
0x16b: frame_vm_group_bin_20000 (RW)
0x16c: frame_vm_group_bin_12801 (RW)
0x16d: frame_vm_group_bin_5736 (RW)
0x16e: frame_vm_group_bin_21837 (RW)
0x16f: frame_vm_group_bin_14662 (RW)
0x170: frame_vm_group_bin_7448 (RW)
0x171: frame_vm_group_bin_0296 (RW)
0x172: frame_vm_group_bin_16477 (RW)
0x173: frame_vm_group_bin_9272 (RW)
0x174: frame_vm_group_bin_2114 (RW)
0x175: frame_vm_group_bin_18209 (RW)
0x176: frame_vm_group_bin_11122 (RW)
0x177: frame_vm_group_bin_3937 (RW)
0x178: frame_vm_group_bin_20033 (RW)
0x179: frame_vm_group_bin_12833 (RW)
0x17: frame_vm_group_bin_10241 (RW)
0x17a: frame_vm_group_bin_5762 (RW)
0x17b: frame_vm_group_bin_21871 (RW)
0x17c: frame_vm_group_bin_14696 (RW)
0x17d: frame_vm_group_bin_7482 (RW)
0x17e: frame_vm_group_bin_23225 (RW)
0x17f: frame_vm_group_bin_16511 (RW)
0x180: frame_vm_group_bin_9301 (RW)
0x181: frame_vm_group_bin_2149 (RW)
0x182: frame_vm_group_bin_18243 (RW)
0x183: frame_vm_group_bin_11155 (RW)
0x184: frame_vm_group_bin_3970 (RW)
0x185: frame_vm_group_bin_20067 (RW)
0x186: frame_vm_group_bin_12867 (RW)
0x187: frame_vm_group_bin_5786 (RW)
0x188: frame_vm_group_bin_21904 (RW)
0x189: frame_vm_group_bin_14729 (RW)
0x18: frame_vm_group_bin_3082 (RW)
0x18a: frame_vm_group_bin_7514 (RW)
0x18b: frame_vm_group_bin_0360 (RW)
0x18c: frame_vm_group_bin_16544 (RW)
0x18d: frame_vm_group_bin_9332 (RW)
0x18e: frame_vm_group_bin_2182 (RW)
0x18f: frame_vm_group_bin_18276 (RW)
0x190: frame_vm_group_bin_11188 (RW)
0x191: frame_vm_group_bin_4003 (RW)
0x192: frame_vm_group_bin_20100 (RW)
0x193: frame_vm_group_bin_12900 (RW)
0x194: frame_vm_group_bin_14977 (RW)
0x195: frame_vm_group_bin_21936 (RW)
0x196: frame_vm_group_bin_14761 (RW)
0x197: frame_vm_group_bin_7546 (RW)
0x198: frame_vm_group_bin_0391 (RW)
0x199: frame_vm_group_bin_16576 (RW)
0x19: frame_vm_group_bin_19150 (RW)
0x19a: frame_vm_group_bin_9366 (RW)
0x19b: frame_vm_group_bin_2212 (RW)
0x19c: frame_vm_group_bin_18310 (RW)
0x19d: frame_vm_group_bin_11222 (RW)
0x19e: frame_vm_group_bin_4037 (RW)
0x19f: frame_vm_group_bin_20133 (RW)
0x1: frame_vm_group_bin_4816 (RW)
0x1a0: frame_vm_group_bin_12933 (RW)
0x1a1: frame_vm_group_bin_5831 (RW)
0x1a2: frame_vm_group_bin_21970 (RW)
0x1a3: frame_vm_group_bin_14794 (RW)
0x1a4: frame_vm_group_bin_7579 (RW)
0x1a5: frame_vm_group_bin_0420 (RW)
0x1a6: frame_vm_group_bin_16609 (RW)
0x1a7: frame_vm_group_bin_9400 (RW)
0x1a8: frame_vm_group_bin_2241 (RW)
0x1a9: frame_vm_group_bin_18343 (RW)
0x1a: frame_vm_group_bin_11988 (RW)
0x1aa: frame_vm_group_bin_11255 (RW)
0x1ab: frame_vm_group_bin_4070 (RW)
0x1ac: frame_vm_group_bin_20165 (RW)
0x1ad: frame_vm_group_bin_12966 (RW)
0x1ae: frame_vm_group_bin_0974 (RW)
0x1af: frame_vm_group_bin_22003 (RW)
0x1b0: frame_vm_group_bin_14827 (RW)
0x1b1: frame_vm_group_bin_7612 (RW)
0x1b2: frame_vm_group_bin_0452 (RW)
0x1b3: frame_vm_group_bin_16642 (RW)
0x1b4: frame_vm_group_bin_9433 (RW)
0x1b5: frame_vm_group_bin_2273 (RW)
0x1b6: frame_vm_group_bin_18376 (RW)
0x1b7: frame_vm_group_bin_11288 (RW)
0x1b8: frame_vm_group_bin_4103 (RW)
0x1b9: frame_vm_group_bin_20197 (RW)
0x1b: frame_vm_group_bin_4883 (RW)
0x1ba: frame_vm_group_bin_13002 (RW)
0x1bb: frame_vm_group_bin_5700 (RW)
0x1bc: frame_vm_group_bin_22031 (RW)
0x1bd: frame_vm_group_bin_14861 (RW)
0x1be: frame_vm_group_bin_7646 (RW)
0x1bf: frame_vm_group_bin_0485 (RW)
0x1c0: frame_vm_group_bin_16676 (RW)
0x1c1: frame_vm_group_bin_9467 (RW)
0x1c2: frame_vm_group_bin_2307 (RW)
0x1c3: frame_vm_group_bin_18408 (RW)
0x1c4: frame_vm_group_bin_11322 (RW)
0x1c5: frame_vm_group_bin_4136 (RW)
0x1c6: frame_vm_group_bin_20231 (RW)
0x1c7: frame_vm_group_bin_13035 (RW)
0x1c8: frame_vm_group_bin_10340 (RW)
0x1c9: frame_vm_group_bin_22052 (RW)
0x1c: frame_vm_group_bin_20976 (RW)
0x1ca: frame_vm_group_bin_14894 (RW)
0x1cb: frame_vm_group_bin_7679 (RW)
0x1cc: frame_vm_group_bin_0518 (RW)
0x1cd: frame_vm_group_bin_16708 (RW)
0x1ce: frame_vm_group_bin_9500 (RW)
0x1cf: frame_vm_group_bin_2340 (RW)
0x1d0: frame_vm_group_bin_18441 (RW)
0x1d1: frame_vm_group_bin_11353 (RW)
0x1d2: frame_vm_group_bin_4168 (RW)
0x1d3: frame_vm_group_bin_20264 (RW)
0x1d4: frame_vm_group_bin_13068 (RW)
0x1d5: frame_vm_group_bin_15002 (RW)
0x1d6: frame_vm_group_bin_22078 (RW)
0x1d7: frame_vm_group_bin_14927 (RW)
0x1d8: frame_vm_group_bin_7712 (RW)
0x1d9: frame_vm_group_bin_0550 (RW)
0x1d: frame_vm_group_bin_13808 (RW)
0x1da: frame_vm_group_bin_16743 (RW)
0x1db: frame_vm_group_bin_9534 (RW)
0x1dc: frame_vm_group_bin_2374 (RW)
0x1dd: frame_vm_group_bin_18473 (RW)
0x1de: frame_vm_group_bin_11386 (RW)
0x1df: frame_vm_group_bin_4201 (RW)
0x1e0: frame_vm_group_bin_20297 (RW)
0x1e1: frame_vm_group_bin_13102 (RW)
0x1e2: frame_vm_group_bin_19623 (RW)
0x1e3: frame_vm_group_bin_22110 (RW)
0x1e4: frame_vm_group_bin_14961 (RW)
0x1e5: frame_vm_group_bin_7745 (RW)
0x1e6: frame_vm_group_bin_0582 (RW)
0x1e7: frame_vm_group_bin_16776 (RW)
0x1e8: frame_vm_group_bin_9567 (RW)
0x1e9: frame_vm_group_bin_2407 (RW)
0x1e: frame_vm_group_bin_6619 (RW)
0x1ea: frame_vm_group_bin_18499 (RW)
0x1eb: frame_vm_group_bin_11418 (RW)
0x1ec: frame_vm_group_bin_4234 (RW)
0x1ed: frame_vm_group_bin_20332 (RW)
0x1ee: frame_vm_group_bin_13135 (RW)
0x1ef: frame_vm_group_bin_5982 (RW)
0x1f0: frame_vm_group_bin_22143 (RW)
0x1f1: frame_vm_group_bin_14994 (RW)
0x1f2: frame_vm_group_bin_7778 (RW)
0x1f3: frame_vm_group_bin_0614 (RW)
0x1f4: frame_vm_group_bin_16809 (RW)
0x1f5: frame_vm_group_bin_9600 (RW)
0x1f6: frame_vm_group_bin_2439 (RW)
0x1f7: frame_vm_group_bin_18525 (RW)
0x1f8: frame_vm_group_bin_11451 (RW)
0x1f9: frame_vm_group_bin_4267 (RW)
0x1f: frame_vm_group_bin_22815 (RW)
0x1fa: frame_vm_group_bin_20366 (RW)
0x1fb: frame_vm_group_bin_13169 (RW)
0x1fc: frame_vm_group_bin_6014 (RW)
0x1fd: frame_vm_group_bin_22177 (RW)
0x1fe: frame_vm_group_bin_15028 (RW)
0x1ff: frame_vm_group_bin_7812 (RW)
0x20: frame_vm_group_bin_15632 (RW)
0x21: frame_vm_group_bin_8442 (RW)
0x22: frame_vm_group_bin_1252 (RW)
0x23: frame_vm_group_bin_17458 (RW)
0x24: frame_vm_group_bin_10275 (RW)
0x25: frame_vm_group_bin_3115 (RW)
0x26: frame_vm_group_bin_19184 (RW)
0x27: frame_vm_group_bin_12019 (RW)
0x28: frame_vm_group_bin_4916 (RW)
0x29: frame_vm_group_bin_21009 (RW)
0x2: frame_vm_group_bin_20920 (RW)
0x2a: frame_vm_group_bin_13837 (RW)
0x2b: frame_vm_group_bin_6652 (RW)
0x2c: frame_vm_group_bin_22848 (RW)
0x2d: frame_vm_group_bin_15665 (RW)
0x2e: frame_vm_group_bin_8475 (RW)
0x2f: frame_vm_group_bin_1283 (RW)
0x30: frame_vm_group_bin_12652 (RW)
0x31: frame_vm_group_bin_10308 (RW)
0x32: frame_vm_group_bin_3148 (RW)
0x33: frame_vm_group_bin_19217 (RW)
0x34: frame_vm_group_bin_12049 (RW)
0x35: frame_vm_group_bin_4947 (RW)
0x36: frame_vm_group_bin_21042 (RW)
0x37: frame_vm_group_bin_13866 (RW)
0x38: frame_vm_group_bin_6685 (RW)
0x39: frame_vm_group_bin_22881 (RW)
0x3: frame_vm_group_bin_13740 (RW)
0x3a: frame_vm_group_bin_15699 (RW)
0x3b: frame_vm_group_bin_8509 (RW)
0x3c: frame_vm_group_bin_1316 (RW)
0x3d: frame_vm_group_bin_17398 (RW)
0x3e: frame_vm_group_bin_10342 (RW)
0x3f: frame_vm_group_bin_3182 (RW)
0x40: frame_vm_group_bin_19251 (RW)
0x41: frame_vm_group_bin_12078 (RW)
0x42: frame_vm_group_bin_4979 (RW)
0x43: frame_vm_group_bin_21077 (RW)
0x44: frame_vm_group_bin_13899 (RW)
0x45: frame_vm_group_bin_6718 (RW)
0x46: frame_vm_group_bin_22915 (RW)
0x47: frame_vm_group_bin_15732 (RW)
0x48: frame_vm_group_bin_8541 (RW)
0x49: frame_vm_group_bin_1349 (RW)
0x4: frame_vm_group_bin_6552 (RW)
0x4a: frame_vm_group_bin_17525 (RW)
0x4b: frame_vm_group_bin_10375 (RW)
0x4c: frame_vm_group_bin_3215 (RW)
0x4d: frame_vm_group_bin_19284 (RW)
0x4e: frame_vm_group_bin_12111 (RW)
0x4f: frame_vm_group_bin_5012 (RW)
0x50: frame_vm_group_bin_21110 (RW)
0x51: frame_vm_group_bin_13932 (RW)
0x52: frame_vm_group_bin_6751 (RW)
0x53: frame_vm_group_bin_22948 (RW)
0x54: frame_vm_group_bin_15765 (RW)
0x55: frame_vm_group_bin_8572 (RW)
0x56: frame_vm_group_bin_1383 (RW)
0x57: frame_vm_group_bin_3406 (RW)
0x58: frame_vm_group_bin_10402 (RW)
0x59: frame_vm_group_bin_3247 (RW)
0x5: frame_vm_group_bin_22748 (RW)
0x5a: frame_vm_group_bin_19318 (RW)
0x5b: frame_vm_group_bin_12144 (RW)
0x5c: frame_vm_group_bin_5046 (RW)
0x5d: frame_vm_group_bin_21143 (RW)
0x5e: frame_vm_group_bin_13966 (RW)
0x5f: frame_vm_group_bin_6784 (RW)
0x60: frame_vm_group_bin_22981 (RW)
0x61: frame_vm_group_bin_15798 (RW)
0x62: frame_vm_group_bin_8605 (RW)
0x63: frame_vm_group_bin_1417 (RW)
0x64: frame_vm_group_bin_8018 (RW)
0x65: frame_vm_group_bin_10431 (RW)
0x66: frame_vm_group_bin_3281 (RW)
0x67: frame_vm_group_bin_19351 (RW)
0x68: frame_vm_group_bin_12174 (RW)
0x69: frame_vm_group_bin_5080 (RW)
0x6: frame_vm_group_bin_15565 (RW)
0x6a: frame_vm_group_bin_21176 (RW)
0x6b: frame_vm_group_bin_13999 (RW)
0x6c: frame_vm_group_bin_6815 (RW)
0x6d: frame_vm_group_bin_23013 (RW)
0x6e: frame_vm_group_bin_15830 (RW)
0x6f: frame_vm_group_bin_8638 (RW)
0x70: frame_vm_group_bin_1450 (RW)
0x71: frame_vm_group_bin_12671 (RW)
0x72: frame_vm_group_bin_10461 (RW)
0x73: frame_vm_group_bin_3314 (RW)
0x74: frame_vm_group_bin_19384 (RW)
0x75: frame_vm_group_bin_6919 (RW)
0x76: frame_vm_group_bin_5113 (RW)
0x77: frame_vm_group_bin_21209 (RW)
0x78: frame_vm_group_bin_14032 (RW)
0x79: frame_vm_group_bin_6843 (RW)
0x7: frame_vm_group_bin_8375 (RW)
0x7a: frame_vm_group_bin_23047 (RW)
0x7b: frame_vm_group_bin_15864 (RW)
0x7c: frame_vm_group_bin_8674 (RW)
0x7d: frame_vm_group_bin_1484 (RW)
0x7e: frame_vm_group_bin_17624 (RW)
0x7f: frame_vm_group_bin_10495 (RW)
0x80: frame_vm_group_bin_3348 (RW)
0x81: frame_vm_group_bin_19417 (RW)
0x82: frame_vm_group_bin_12236 (RW)
0x83: frame_vm_group_bin_5147 (RW)
0x84: frame_vm_group_bin_21243 (RW)
0x85: frame_vm_group_bin_14066 (RW)
0x86: frame_vm_group_bin_6872 (RW)
0x87: frame_vm_group_bin_23080 (RW)
0x88: frame_vm_group_bin_15897 (RW)
0x89: frame_vm_group_bin_8706 (RW)
0x8: frame_vm_group_bin_1186 (RW)
0x8a: frame_vm_group_bin_1517 (RW)
0x8b: frame_vm_group_bin_17657 (RW)
0x8c: frame_vm_group_bin_10527 (RW)
0x8d: frame_vm_group_bin_3379 (RW)
0x8e: frame_vm_group_bin_19448 (RW)
0x8f: frame_vm_group_bin_12269 (RW)
0x90: frame_vm_group_bin_5180 (RW)
0x91: frame_vm_group_bin_21276 (RW)
0x92: frame_vm_group_bin_14099 (RW)
0x93: frame_vm_group_bin_6895 (RW)
0x94: frame_vm_group_bin_23113 (RW)
0x95: frame_vm_group_bin_15930 (RW)
0x96: frame_vm_group_bin_8739 (RW)
0x97: frame_vm_group_bin_1550 (RW)
0x98: frame_vm_group_bin_3425 (RW)
0x99: frame_vm_group_bin_10560 (RW)
0x9: frame_vm_group_bin_17406 (RW)
0x9a: frame_vm_group_bin_3407 (RW)
0x9b: frame_vm_group_bin_19481 (RW)
0x9c: frame_vm_group_bin_12303 (RW)
0x9d: frame_vm_group_bin_5214 (RW)
0x9e: frame_vm_group_bin_21309 (RW)
0x9f: frame_vm_group_bin_14133 (RW)
0xa0: frame_vm_group_bin_6923 (RW)
0xa1: frame_vm_group_bin_23146 (RW)
0xa2: frame_vm_group_bin_15964 (RW)
0xa3: frame_vm_group_bin_8773 (RW)
0xa4: frame_vm_group_bin_1584 (RW)
0xa5: frame_vm_group_bin_8037 (RW)
0xa6: frame_vm_group_bin_10594 (RW)
0xa7: frame_vm_group_bin_3432 (RW)
0xa8: frame_vm_group_bin_19514 (RW)
0xa9: frame_vm_group_bin_12335 (RW)
0xa: frame_vm_group_bin_10208 (RW)
0xaa: frame_vm_group_bin_5247 (RW)
0xab: frame_vm_group_bin_21341 (RW)
0xac: frame_vm_group_bin_14166 (RW)
0xad: frame_vm_group_bin_6953 (RW)
0xae: frame_vm_group_bin_23179 (RW)
0xaf: frame_vm_group_bin_15999 (RW)
0xb0: frame_vm_group_bin_8806 (RW)
0xb1: frame_vm_group_bin_1617 (RW)
0xb2: frame_vm_group_bin_12687 (RW)
0xb3: frame_vm_group_bin_10627 (RW)
0xb4: frame_vm_group_bin_3454 (RW)
0xb5: frame_vm_group_bin_19547 (RW)
0xb6: frame_vm_group_bin_12368 (RW)
0xb7: frame_vm_group_bin_5280 (RW)
0xb8: frame_vm_group_bin_21374 (RW)
0xb9: frame_vm_group_bin_14198 (RW)
0xb: frame_vm_group_bin_3049 (RW)
0xba: frame_vm_group_bin_6986 (RW)
0xbb: frame_vm_group_bin_23209 (RW)
0xbc: frame_vm_group_bin_16033 (RW)
0xbd: frame_vm_group_bin_8840 (RW)
0xbe: frame_vm_group_bin_1651 (RW)
0xbf: frame_vm_group_bin_17434 (RW)
0xc0: frame_vm_group_bin_10659 (RW)
0xc1: frame_vm_group_bin_3483 (RW)
0xc2: frame_vm_group_bin_19582 (RW)
0xc3: frame_vm_group_bin_12402 (RW)
0xc4: frame_vm_group_bin_5313 (RW)
0xc5: frame_vm_group_bin_21408 (RW)
0xc6: frame_vm_group_bin_14232 (RW)
0xc7: frame_vm_group_bin_7019 (RW)
0xc8: frame_vm_group_bin_23231 (RW)
0xc9: frame_vm_group_bin_16066 (RW)
0xc: frame_vm_group_bin_19118 (RW)
0xca: frame_vm_group_bin_8872 (RW)
0xcb: frame_vm_group_bin_1684 (RW)
0xcc: frame_vm_group_bin_17801 (RW)
0xcd: frame_vm_group_bin_10692 (RW)
0xce: frame_vm_group_bin_3509 (RW)
0xcf: frame_vm_group_bin_19615 (RW)
0xd0: frame_vm_group_bin_12434 (RW)
0xd1: frame_vm_group_bin_5345 (RW)
0xd2: frame_vm_group_bin_21440 (RW)
0xd3: frame_vm_group_bin_14264 (RW)
0xd4: frame_vm_group_bin_7051 (RW)
0xd5: frame_vm_group_bin_23252 (RW)
0xd6: frame_vm_group_bin_16098 (RW)
0xd7: frame_vm_group_bin_8904 (RW)
0xd8: frame_vm_group_bin_1716 (RW)
0xd9: frame_vm_group_bin_3440 (RW)
0xd: frame_vm_group_bin_11954 (RW)
0xda: frame_vm_group_bin_10725 (RW)
0xdb: frame_vm_group_bin_3539 (RW)
0xdc: frame_vm_group_bin_19647 (RW)
0xdd: frame_vm_group_bin_12467 (RW)
0xde: frame_vm_group_bin_5377 (RW)
0xdf: frame_vm_group_bin_21473 (RW)
0xe0: frame_vm_group_bin_14296 (RW)
0xe1: frame_vm_group_bin_7083 (RW)
0xe2: frame_vm_group_bin_13807 (RW)
0xe3: frame_vm_group_bin_16130 (RW)
0xe4: frame_vm_group_bin_8937 (RW)
0xe5: frame_vm_group_bin_1749 (RW)
0xe6: frame_vm_group_bin_17858 (RW)
0xe7: frame_vm_group_bin_10757 (RW)
0xe8: frame_vm_group_bin_3570 (RW)
0xe9: frame_vm_group_bin_19674 (RW)
0xe: frame_vm_group_bin_4849 (RW)
0xea: frame_vm_group_bin_12499 (RW)
0xeb: frame_vm_group_bin_5409 (RW)
0xec: frame_vm_group_bin_21504 (RW)
0xed: frame_vm_group_bin_14328 (RW)
0xee: frame_vm_group_bin_7114 (RW)
0xef: frame_vm_group_bin_0039 (RW)
0xf0: frame_vm_group_bin_16162 (RW)
0xf1: frame_vm_group_bin_8969 (RW)
0xf2: frame_vm_group_bin_1781 (RW)
0xf3: frame_vm_group_bin_17885 (RW)
0xf4: frame_vm_group_bin_10789 (RW)
0xf5: frame_vm_group_bin_3604 (RW)
0xf6: frame_vm_group_bin_19704 (RW)
0xf7: frame_vm_group_bin_12532 (RW)
0xf8: frame_vm_group_bin_5442 (RW)
0xf9: frame_vm_group_bin_21537 (RW)
0xf: frame_vm_group_bin_20947 (RW)
0xfa: frame_vm_group_bin_14362 (RW)
0xfb: frame_vm_group_bin_7147 (RW)
0xfc: frame_vm_group_bin_0065 (RW)
0xfd: frame_vm_group_bin_16196 (RW)
0xfe: frame_vm_group_bin_9003 (RW)
0xff: frame_vm_group_bin_1815 (RW)
}
pt_vm_group_bin_0065 {
0x0: frame_vm_group_bin_6455 (RW)
0x100: frame_vm_group_bin_12470 (RW)
0x101: frame_vm_group_bin_5380 (RW)
0x102: frame_vm_group_bin_21476 (RW)
0x103: frame_vm_group_bin_14299 (RW)
0x104: frame_vm_group_bin_7086 (RW)
0x105: frame_vm_group_bin_21918 (RW)
0x106: frame_vm_group_bin_16133 (RW)
0x107: frame_vm_group_bin_8940 (RW)
0x108: frame_vm_group_bin_1752 (RW)
0x109: frame_vm_group_bin_17860 (RW)
0x10: frame_vm_group_bin_8311 (RW)
0x10a: frame_vm_group_bin_10760 (RW)
0x10b: frame_vm_group_bin_3573 (RW)
0x10c: frame_vm_group_bin_11843 (RW)
0x10d: frame_vm_group_bin_12502 (RW)
0x10e: frame_vm_group_bin_5412 (RW)
0x10f: frame_vm_group_bin_21507 (RW)
0x110: frame_vm_group_bin_14331 (RW)
0x111: frame_vm_group_bin_7117 (RW)
0x112: frame_vm_group_bin_0040 (RW)
0x113: frame_vm_group_bin_16165 (RW)
0x114: frame_vm_group_bin_8972 (RW)
0x115: frame_vm_group_bin_1784 (RW)
0x116: frame_vm_group_bin_17888 (RW)
0x117: frame_vm_group_bin_10792 (RW)
0x118: frame_vm_group_bin_3607 (RW)
0x119: frame_vm_group_bin_19707 (RW)
0x11: frame_vm_group_bin_1122 (RW)
0x11a: frame_vm_group_bin_12536 (RW)
0x11b: frame_vm_group_bin_5446 (RW)
0x11c: frame_vm_group_bin_21541 (RW)
0x11d: frame_vm_group_bin_14365 (RW)
0x11e: frame_vm_group_bin_7150 (RW)
0x11f: frame_vm_group_bin_7902 (RW)
0x120: frame_vm_group_bin_16199 (RW)
0x121: frame_vm_group_bin_9006 (RW)
0x122: frame_vm_group_bin_1818 (RW)
0x123: frame_vm_group_bin_17920 (RW)
0x124: frame_vm_group_bin_10826 (RW)
0x125: frame_vm_group_bin_3641 (RW)
0x126: frame_vm_group_bin_19741 (RW)
0x127: frame_vm_group_bin_12569 (RW)
0x128: frame_vm_group_bin_5477 (RW)
0x129: frame_vm_group_bin_21574 (RW)
0x12: frame_vm_group_bin_17348 (RW)
0x12a: frame_vm_group_bin_14398 (RW)
0x12b: frame_vm_group_bin_7185 (RW)
0x12c: frame_vm_group_bin_0092 (RW)
0x12d: frame_vm_group_bin_16226 (RW)
0x12e: frame_vm_group_bin_9039 (RW)
0x12f: frame_vm_group_bin_1851 (RW)
0x130: frame_vm_group_bin_17951 (RW)
0x131: frame_vm_group_bin_10859 (RW)
0x132: frame_vm_group_bin_3674 (RW)
0x133: frame_vm_group_bin_19774 (RW)
0x134: frame_vm_group_bin_12602 (RW)
0x135: frame_vm_group_bin_5510 (RW)
0x136: frame_vm_group_bin_21607 (RW)
0x137: frame_vm_group_bin_14431 (RW)
0x138: frame_vm_group_bin_7218 (RW)
0x139: frame_vm_group_bin_0117 (RW)
0x13: frame_vm_group_bin_10142 (RW)
0x13a: frame_vm_group_bin_16253 (RW)
0x13b: frame_vm_group_bin_9073 (RW)
0x13c: frame_vm_group_bin_1885 (RW)
0x13d: frame_vm_group_bin_17983 (RW)
0x13e: frame_vm_group_bin_10893 (RW)
0x13f: frame_vm_group_bin_3708 (RW)
0x140: frame_vm_group_bin_19808 (RW)
0x141: frame_vm_group_bin_12636 (RW)
0x142: frame_vm_group_bin_5543 (RW)
0x143: frame_vm_group_bin_21641 (RW)
0x144: frame_vm_group_bin_14465 (RW)
0x145: frame_vm_group_bin_7252 (RW)
0x146: frame_vm_group_bin_0139 (RW)
0x147: frame_vm_group_bin_20484 (RW)
0x148: frame_vm_group_bin_9106 (RW)
0x149: frame_vm_group_bin_1918 (RW)
0x14: frame_vm_group_bin_2985 (RW)
0x14a: frame_vm_group_bin_18016 (RW)
0x14b: frame_vm_group_bin_10926 (RW)
0x14c: frame_vm_group_bin_3741 (RW)
0x14d: frame_vm_group_bin_19841 (RW)
0x14e: frame_vm_group_bin_12665 (RW)
0x14f: frame_vm_group_bin_5576 (RW)
0x150: frame_vm_group_bin_21674 (RW)
0x151: frame_vm_group_bin_14498 (RW)
0x152: frame_vm_group_bin_7285 (RW)
0x153: frame_vm_group_bin_0161 (RW)
0x154: frame_vm_group_bin_16314 (RW)
0x155: frame_vm_group_bin_9139 (RW)
0x156: frame_vm_group_bin_1951 (RW)
0x157: frame_vm_group_bin_18049 (RW)
0x158: frame_vm_group_bin_10959 (RW)
0x159: frame_vm_group_bin_3774 (RW)
0x15: frame_vm_group_bin_19055 (RW)
0x15a: frame_vm_group_bin_19875 (RW)
0x15b: frame_vm_group_bin_12689 (RW)
0x15c: frame_vm_group_bin_5609 (RW)
0x15d: frame_vm_group_bin_21707 (RW)
0x15e: frame_vm_group_bin_14533 (RW)
0x15f: frame_vm_group_bin_7318 (RW)
0x160: frame_vm_group_bin_0192 (RW)
0x161: frame_vm_group_bin_16347 (RW)
0x162: frame_vm_group_bin_9171 (RW)
0x163: frame_vm_group_bin_1984 (RW)
0x164: frame_vm_group_bin_18081 (RW)
0x165: frame_vm_group_bin_10992 (RW)
0x166: frame_vm_group_bin_3807 (RW)
0x167: frame_vm_group_bin_19906 (RW)
0x168: frame_vm_group_bin_19754 (RW)
0x169: frame_vm_group_bin_5640 (RW)
0x16: frame_vm_group_bin_11897 (RW)
0x16a: frame_vm_group_bin_21740 (RW)
0x16b: frame_vm_group_bin_14566 (RW)
0x16c: frame_vm_group_bin_7351 (RW)
0x16d: frame_vm_group_bin_0223 (RW)
0x16e: frame_vm_group_bin_16380 (RW)
0x16f: frame_vm_group_bin_9202 (RW)
0x170: frame_vm_group_bin_2017 (RW)
0x171: frame_vm_group_bin_18113 (RW)
0x172: frame_vm_group_bin_11025 (RW)
0x173: frame_vm_group_bin_3840 (RW)
0x174: frame_vm_group_bin_19938 (RW)
0x175: frame_vm_group_bin_1105 (RW)
0x176: frame_vm_group_bin_5673 (RW)
0x177: frame_vm_group_bin_21773 (RW)
0x178: frame_vm_group_bin_14599 (RW)
0x179: frame_vm_group_bin_7384 (RW)
0x17: frame_vm_group_bin_4786 (RW)
0x17a: frame_vm_group_bin_0247 (RW)
0x17b: frame_vm_group_bin_16414 (RW)
0x17c: frame_vm_group_bin_14411 (RW)
0x17d: frame_vm_group_bin_2051 (RW)
0x17e: frame_vm_group_bin_18147 (RW)
0x17f: frame_vm_group_bin_11059 (RW)
0x180: frame_vm_group_bin_3874 (RW)
0x181: frame_vm_group_bin_19972 (RW)
0x182: frame_vm_group_bin_12771 (RW)
0x183: frame_vm_group_bin_5707 (RW)
0x184: frame_vm_group_bin_21807 (RW)
0x185: frame_vm_group_bin_14632 (RW)
0x186: frame_vm_group_bin_7418 (RW)
0x187: frame_vm_group_bin_0270 (RW)
0x188: frame_vm_group_bin_16447 (RW)
0x189: frame_vm_group_bin_19035 (RW)
0x18: frame_vm_group_bin_20894 (RW)
0x18a: frame_vm_group_bin_2084 (RW)
0x18b: frame_vm_group_bin_18180 (RW)
0x18c: frame_vm_group_bin_11092 (RW)
0x18d: frame_vm_group_bin_3907 (RW)
0x18e: frame_vm_group_bin_20003 (RW)
0x18f: frame_vm_group_bin_12804 (RW)
0x190: frame_vm_group_bin_5739 (RW)
0x191: frame_vm_group_bin_21840 (RW)
0x192: frame_vm_group_bin_14665 (RW)
0x193: frame_vm_group_bin_7451 (RW)
0x194: frame_vm_group_bin_0299 (RW)
0x195: frame_vm_group_bin_16480 (RW)
0x196: frame_vm_group_bin_9275 (RW)
0x197: frame_vm_group_bin_2117 (RW)
0x198: frame_vm_group_bin_18212 (RW)
0x199: frame_vm_group_bin_19413 (RW)
0x19: frame_vm_group_bin_13710 (RW)
0x19a: frame_vm_group_bin_20316 (RW)
0x19b: frame_vm_group_bin_20037 (RW)
0x19c: frame_vm_group_bin_12837 (RW)
0x19d: frame_vm_group_bin_13687 (RW)
0x19e: frame_vm_group_bin_21874 (RW)
0x19f: frame_vm_group_bin_14699 (RW)
0x1: frame_vm_group_bin_22652 (RW)
0x1a0: frame_vm_group_bin_7485 (RW)
0x1a1: frame_vm_group_bin_0331 (RW)
0x1a2: frame_vm_group_bin_16514 (RW)
0x1a3: frame_vm_group_bin_9304 (RW)
0x1a4: frame_vm_group_bin_2152 (RW)
0x1a5: frame_vm_group_bin_18246 (RW)
0x1a6: frame_vm_group_bin_11158 (RW)
0x1a7: frame_vm_group_bin_3973 (RW)
0x1a8: frame_vm_group_bin_20070 (RW)
0x1a9: frame_vm_group_bin_12870 (RW)
0x1a: frame_vm_group_bin_6522 (RW)
0x1aa: frame_vm_group_bin_18333 (RW)
0x1ab: frame_vm_group_bin_21907 (RW)
0x1ac: frame_vm_group_bin_14732 (RW)
0x1ad: frame_vm_group_bin_7517 (RW)
0x1ae: frame_vm_group_bin_0363 (RW)
0x1af: frame_vm_group_bin_16547 (RW)
0x1b0: frame_vm_group_bin_9335 (RW)
0x1b1: frame_vm_group_bin_2185 (RW)
0x1b2: frame_vm_group_bin_18279 (RW)
0x1b3: frame_vm_group_bin_11191 (RW)
0x1b4: frame_vm_group_bin_4006 (RW)
0x1b5: frame_vm_group_bin_20103 (RW)
0x1b6: frame_vm_group_bin_12903 (RW)
0x1b7: frame_vm_group_bin_23071 (RW)
0x1b8: frame_vm_group_bin_21939 (RW)
0x1b9: frame_vm_group_bin_14764 (RW)
0x1b: frame_vm_group_bin_22719 (RW)
0x1ba: frame_vm_group_bin_18683 (RW)
0x1bb: frame_vm_group_bin_0395 (RW)
0x1bc: frame_vm_group_bin_16580 (RW)
0x1bd: frame_vm_group_bin_9369 (RW)
0x1be: frame_vm_group_bin_2215 (RW)
0x1bf: frame_vm_group_bin_18313 (RW)
0x1c0: frame_vm_group_bin_11225 (RW)
0x1c1: frame_vm_group_bin_4040 (RW)
0x1c2: frame_vm_group_bin_20136 (RW)
0x1c3: frame_vm_group_bin_12936 (RW)
0x1c4: frame_vm_group_bin_5832 (RW)
0x1c5: frame_vm_group_bin_21973 (RW)
0x1c6: frame_vm_group_bin_14797 (RW)
0x1c7: frame_vm_group_bin_7582 (RW)
0x1c8: frame_vm_group_bin_0422 (RW)
0x1c9: frame_vm_group_bin_16612 (RW)
0x1c: frame_vm_group_bin_15536 (RW)
0x1ca: frame_vm_group_bin_9403 (RW)
0x1cb: frame_vm_group_bin_17645 (RW)
0x1cc: frame_vm_group_bin_18346 (RW)
0x1cd: frame_vm_group_bin_11258 (RW)
0x1ce: frame_vm_group_bin_4073 (RW)
0x1cf: frame_vm_group_bin_20168 (RW)
0x1d0: frame_vm_group_bin_12969 (RW)
0x1d1: frame_vm_group_bin_5856 (RW)
0x1d2: frame_vm_group_bin_22006 (RW)
0x1d3: frame_vm_group_bin_14830 (RW)
0x1d4: frame_vm_group_bin_7615 (RW)
0x1d5: frame_vm_group_bin_0455 (RW)
0x1d6: frame_vm_group_bin_16645 (RW)
0x1d7: frame_vm_group_bin_9436 (RW)
0x1d8: frame_vm_group_bin_2276 (RW)
0x1d9: frame_vm_group_bin_18379 (RW)
0x1d: frame_vm_group_bin_8345 (RW)
0x1da: frame_vm_group_bin_11292 (RW)
0x1db: frame_vm_group_bin_4107 (RW)
0x1dc: frame_vm_group_bin_20201 (RW)
0x1dd: frame_vm_group_bin_13005 (RW)
0x1de: frame_vm_group_bin_5882 (RW)
0x1df: frame_vm_group_bin_22034 (RW)
0x1e0: frame_vm_group_bin_14864 (RW)
0x1e1: frame_vm_group_bin_7649 (RW)
0x1e2: frame_vm_group_bin_0488 (RW)
0x1e3: frame_vm_group_bin_16679 (RW)
0x1e4: frame_vm_group_bin_9470 (RW)
0x1e5: frame_vm_group_bin_2310 (RW)
0x1e6: frame_vm_group_bin_18411 (RW)
0x1e7: frame_vm_group_bin_11325 (RW)
0x1e8: frame_vm_group_bin_4139 (RW)
0x1e9: frame_vm_group_bin_20234 (RW)
0x1e: frame_vm_group_bin_1156 (RW)
0x1ea: frame_vm_group_bin_13038 (RW)
0x1eb: frame_vm_group_bin_5908 (RW)
0x1ec: frame_vm_group_bin_17002 (RW)
0x1ed: frame_vm_group_bin_14897 (RW)
0x1ee: frame_vm_group_bin_7682 (RW)
0x1ef: frame_vm_group_bin_0521 (RW)
0x1f0: frame_vm_group_bin_16711 (RW)
0x1f1: frame_vm_group_bin_9503 (RW)
0x1f2: frame_vm_group_bin_2343 (RW)
0x1f3: frame_vm_group_bin_18444 (RW)
0x1f4: frame_vm_group_bin_11356 (RW)
0x1f5: frame_vm_group_bin_4171 (RW)
0x1f6: frame_vm_group_bin_20267 (RW)
0x1f7: frame_vm_group_bin_13071 (RW)
0x1f8: frame_vm_group_bin_5933 (RW)
0x1f9: frame_vm_group_bin_22081 (RW)
0x1f: frame_vm_group_bin_17381 (RW)
0x1fa: frame_vm_group_bin_14931 (RW)
0x1fb: frame_vm_group_bin_7716 (RW)
0x1fc: frame_vm_group_bin_0553 (RW)
0x1fd: frame_vm_group_bin_16746 (RW)
0x1fe: frame_vm_group_bin_9537 (RW)
0x1ff: frame_vm_group_bin_2377 (RW)
0x20: frame_vm_group_bin_10178 (RW)
0x21: frame_vm_group_bin_3019 (RW)
0x22: frame_vm_group_bin_19089 (RW)
0x23: frame_vm_group_bin_11927 (RW)
0x24: frame_vm_group_bin_4819 (RW)
0x25: frame_vm_group_bin_16838 (RW)
0x26: frame_vm_group_bin_13743 (RW)
0x27: frame_vm_group_bin_6555 (RW)
0x28: frame_vm_group_bin_22751 (RW)
0x29: frame_vm_group_bin_15568 (RW)
0x2: frame_vm_group_bin_15470 (RW)
0x2a: frame_vm_group_bin_8378 (RW)
0x2b: frame_vm_group_bin_1189 (RW)
0x2c: frame_vm_group_bin_17409 (RW)
0x2d: frame_vm_group_bin_10211 (RW)
0x2e: frame_vm_group_bin_3052 (RW)
0x2f: frame_vm_group_bin_19121 (RW)
0x30: frame_vm_group_bin_11957 (RW)
0x31: frame_vm_group_bin_4852 (RW)
0x32: frame_vm_group_bin_21470 (RW)
0x33: frame_vm_group_bin_13777 (RW)
0x34: frame_vm_group_bin_6588 (RW)
0x35: frame_vm_group_bin_22784 (RW)
0x36: frame_vm_group_bin_15601 (RW)
0x37: frame_vm_group_bin_8411 (RW)
0x38: frame_vm_group_bin_1222 (RW)
0x39: frame_vm_group_bin_17433 (RW)
0x3: frame_vm_group_bin_8278 (RW)
0x3a: frame_vm_group_bin_10245 (RW)
0x3b: frame_vm_group_bin_3086 (RW)
0x3c: frame_vm_group_bin_19154 (RW)
0x3d: frame_vm_group_bin_5744 (RW)
0x3e: frame_vm_group_bin_4886 (RW)
0x3f: frame_vm_group_bin_20979 (RW)
0x40: frame_vm_group_bin_13811 (RW)
0x41: frame_vm_group_bin_6622 (RW)
0x42: frame_vm_group_bin_22818 (RW)
0x43: frame_vm_group_bin_15635 (RW)
0x44: frame_vm_group_bin_8445 (RW)
0x45: frame_vm_group_bin_1255 (RW)
0x46: frame_vm_group_bin_16124 (RW)
0x47: frame_vm_group_bin_10278 (RW)
0x48: frame_vm_group_bin_3118 (RW)
0x49: frame_vm_group_bin_19187 (RW)
0x4: frame_vm_group_bin_17516 (RW)
0x4a: frame_vm_group_bin_12021 (RW)
0x4b: frame_vm_group_bin_4919 (RW)
0x4c: frame_vm_group_bin_21012 (RW)
0x4d: frame_vm_group_bin_13840 (RW)
0x4e: frame_vm_group_bin_6655 (RW)
0x4f: frame_vm_group_bin_22851 (RW)
0x50: frame_vm_group_bin_15668 (RW)
0x51: frame_vm_group_bin_8478 (RW)
0x52: frame_vm_group_bin_1286 (RW)
0x53: frame_vm_group_bin_17476 (RW)
0x54: frame_vm_group_bin_10311 (RW)
0x55: frame_vm_group_bin_3151 (RW)
0x56: frame_vm_group_bin_19220 (RW)
0x57: frame_vm_group_bin_12050 (RW)
0x58: frame_vm_group_bin_4950 (RW)
0x59: frame_vm_group_bin_21046 (RW)
0x5: frame_vm_group_bin_17315 (RW)
0x5a: frame_vm_group_bin_13870 (RW)
0x5b: frame_vm_group_bin_6689 (RW)
0x5c: frame_vm_group_bin_22885 (RW)
0x5d: frame_vm_group_bin_15702 (RW)
0x5e: frame_vm_group_bin_5020 (RW)
0x5f: frame_vm_group_bin_1319 (RW)
0x60: frame_vm_group_bin_2121 (RW)
0x61: frame_vm_group_bin_10345 (RW)
0x62: frame_vm_group_bin_3185 (RW)
0x63: frame_vm_group_bin_19254 (RW)
0x64: frame_vm_group_bin_12081 (RW)
0x65: frame_vm_group_bin_4982 (RW)
0x66: frame_vm_group_bin_21080 (RW)
0x67: frame_vm_group_bin_13902 (RW)
0x68: frame_vm_group_bin_6721 (RW)
0x69: frame_vm_group_bin_22918 (RW)
0x6: frame_vm_group_bin_10109 (RW)
0x6a: frame_vm_group_bin_15735 (RW)
0x6b: frame_vm_group_bin_8544 (RW)
0x6c: frame_vm_group_bin_1352 (RW)
0x6d: frame_vm_group_bin_17527 (RW)
0x6e: frame_vm_group_bin_10378 (RW)
0x6f: frame_vm_group_bin_3218 (RW)
0x70: frame_vm_group_bin_19287 (RW)
0x71: frame_vm_group_bin_12113 (RW)
0x72: frame_vm_group_bin_5015 (RW)
0x73: frame_vm_group_bin_21113 (RW)
0x74: frame_vm_group_bin_13935 (RW)
0x75: frame_vm_group_bin_6754 (RW)
0x76: frame_vm_group_bin_22951 (RW)
0x77: frame_vm_group_bin_15768 (RW)
0x78: frame_vm_group_bin_8575 (RW)
0x79: frame_vm_group_bin_1386 (RW)
0x7: frame_vm_group_bin_2952 (RW)
0x7a: frame_vm_group_bin_17552 (RW)
0x7b: frame_vm_group_bin_10029 (RW)
0x7c: frame_vm_group_bin_3251 (RW)
0x7d: frame_vm_group_bin_19321 (RW)
0x7e: frame_vm_group_bin_12147 (RW)
0x7f: frame_vm_group_bin_5049 (RW)
0x80: frame_vm_group_bin_21146 (RW)
0x81: frame_vm_group_bin_13969 (RW)
0x82: frame_vm_group_bin_6787 (RW)
0x83: frame_vm_group_bin_22984 (RW)
0x84: frame_vm_group_bin_15801 (RW)
0x85: frame_vm_group_bin_8608 (RW)
0x86: frame_vm_group_bin_1420 (RW)
0x87: frame_vm_group_bin_17573 (RW)
0x88: frame_vm_group_bin_10434 (RW)
0x89: frame_vm_group_bin_3284 (RW)
0x8: frame_vm_group_bin_19022 (RW)
0x8a: frame_vm_group_bin_19354 (RW)
0x8b: frame_vm_group_bin_12177 (RW)
0x8c: frame_vm_group_bin_5083 (RW)
0x8d: frame_vm_group_bin_21179 (RW)
0x8e: frame_vm_group_bin_14002 (RW)
0x8f: frame_vm_group_bin_6818 (RW)
0x90: frame_vm_group_bin_23016 (RW)
0x91: frame_vm_group_bin_15833 (RW)
0x92: frame_vm_group_bin_8641 (RW)
0x93: frame_vm_group_bin_1453 (RW)
0x94: frame_vm_group_bin_17596 (RW)
0x95: frame_vm_group_bin_10464 (RW)
0x96: frame_vm_group_bin_3317 (RW)
0x97: frame_vm_group_bin_19387 (RW)
0x98: frame_vm_group_bin_15062 (RW)
0x99: frame_vm_group_bin_5116 (RW)
0x9: frame_vm_group_bin_11874 (RW)
0x9a: frame_vm_group_bin_21213 (RW)
0x9b: frame_vm_group_bin_14036 (RW)
0x9c: frame_vm_group_bin_6847 (RW)
0x9d: frame_vm_group_bin_23050 (RW)
0x9e: frame_vm_group_bin_15867 (RW)
0x9f: frame_vm_group_bin_8677 (RW)
0xa0: frame_vm_group_bin_1487 (RW)
0xa1: frame_vm_group_bin_17627 (RW)
0xa2: frame_vm_group_bin_10498 (RW)
0xa3: frame_vm_group_bin_3351 (RW)
0xa4: frame_vm_group_bin_19420 (RW)
0xa5: frame_vm_group_bin_12239 (RW)
0xa6: frame_vm_group_bin_5150 (RW)
0xa7: frame_vm_group_bin_21246 (RW)
0xa8: frame_vm_group_bin_14069 (RW)
0xa9: frame_vm_group_bin_13964 (RW)
0xa: frame_vm_group_bin_4753 (RW)
0xaa: frame_vm_group_bin_23083 (RW)
0xab: frame_vm_group_bin_15900 (RW)
0xac: frame_vm_group_bin_8709 (RW)
0xad: frame_vm_group_bin_1520 (RW)
0xae: frame_vm_group_bin_17660 (RW)
0xaf: frame_vm_group_bin_10530 (RW)
0xb0: frame_vm_group_bin_3382 (RW)
0xb1: frame_vm_group_bin_19451 (RW)
0xb2: frame_vm_group_bin_12272 (RW)
0xb3: frame_vm_group_bin_5183 (RW)
0xb4: frame_vm_group_bin_21279 (RW)
0xb5: frame_vm_group_bin_14102 (RW)
0xb6: frame_vm_group_bin_18590 (RW)
0xb7: frame_vm_group_bin_23116 (RW)
0xb8: frame_vm_group_bin_15933 (RW)
0xb9: frame_vm_group_bin_8742 (RW)
0xb: frame_vm_group_bin_20868 (RW)
0xba: frame_vm_group_bin_1554 (RW)
0xbb: frame_vm_group_bin_17690 (RW)
0xbc: frame_vm_group_bin_10564 (RW)
0xbd: frame_vm_group_bin_3410 (RW)
0xbe: frame_vm_group_bin_19484 (RW)
0xbf: frame_vm_group_bin_12306 (RW)
0xc0: frame_vm_group_bin_5217 (RW)
0xc1: frame_vm_group_bin_21312 (RW)
0xc2: frame_vm_group_bin_14136 (RW)
0xc3: frame_vm_group_bin_6926 (RW)
0xc4: frame_vm_group_bin_23149 (RW)
0xc5: frame_vm_group_bin_15967 (RW)
0xc6: frame_vm_group_bin_8776 (RW)
0xc7: frame_vm_group_bin_1587 (RW)
0xc8: frame_vm_group_bin_17716 (RW)
0xc9: frame_vm_group_bin_10597 (RW)
0xc: frame_vm_group_bin_13677 (RW)
0xca: frame_vm_group_bin_13240 (RW)
0xcb: frame_vm_group_bin_19517 (RW)
0xcc: frame_vm_group_bin_12338 (RW)
0xcd: frame_vm_group_bin_5250 (RW)
0xce: frame_vm_group_bin_21344 (RW)
0xcf: frame_vm_group_bin_14169 (RW)
0xd0: frame_vm_group_bin_6956 (RW)
0xd1: frame_vm_group_bin_23182 (RW)
0xd2: frame_vm_group_bin_16002 (RW)
0xd3: frame_vm_group_bin_8809 (RW)
0xd4: frame_vm_group_bin_1620 (RW)
0xd5: frame_vm_group_bin_17742 (RW)
0xd6: frame_vm_group_bin_10630 (RW)
0xd7: frame_vm_group_bin_17892 (RW)
0xd8: frame_vm_group_bin_19550 (RW)
0xd9: frame_vm_group_bin_12371 (RW)
0xd: frame_vm_group_bin_6488 (RW)
0xda: frame_vm_group_bin_5284 (RW)
0xdb: frame_vm_group_bin_21378 (RW)
0xdc: frame_vm_group_bin_14202 (RW)
0xdd: frame_vm_group_bin_6989 (RW)
0xde: frame_vm_group_bin_23212 (RW)
0xdf: frame_vm_group_bin_16036 (RW)
0xe0: frame_vm_group_bin_8843 (RW)
0xe1: frame_vm_group_bin_1654 (RW)
0xe2: frame_vm_group_bin_17773 (RW)
0xe3: frame_vm_group_bin_10662 (RW)
0xe4: frame_vm_group_bin_22623 (RW)
0xe5: frame_vm_group_bin_19585 (RW)
0xe6: frame_vm_group_bin_12405 (RW)
0xe7: frame_vm_group_bin_5316 (RW)
0xe8: frame_vm_group_bin_21411 (RW)
0xe9: frame_vm_group_bin_14235 (RW)
0xe: frame_vm_group_bin_22685 (RW)
0xea: frame_vm_group_bin_7022 (RW)
0xeb: frame_vm_group_bin_12535 (RW)
0xec: frame_vm_group_bin_16069 (RW)
0xed: frame_vm_group_bin_8875 (RW)
0xee: frame_vm_group_bin_1687 (RW)
0xef: frame_vm_group_bin_17804 (RW)
0xf0: frame_vm_group_bin_10695 (RW)
0xf1: frame_vm_group_bin_3986 (RW)
0xf2: frame_vm_group_bin_19618 (RW)
0xf3: frame_vm_group_bin_12437 (RW)
0xf4: frame_vm_group_bin_5348 (RW)
0xf5: frame_vm_group_bin_21443 (RW)
0xf6: frame_vm_group_bin_14267 (RW)
0xf7: frame_vm_group_bin_7054 (RW)
0xf8: frame_vm_group_bin_23255 (RW)
0xf9: frame_vm_group_bin_16101 (RW)
0xf: frame_vm_group_bin_15503 (RW)
0xfa: frame_vm_group_bin_8908 (RW)
0xfb: frame_vm_group_bin_1720 (RW)
0xfc: frame_vm_group_bin_17833 (RW)
0xfd: frame_vm_group_bin_10728 (RW)
0xfe: frame_vm_group_bin_3542 (RW)
0xff: frame_vm_group_bin_19650 (RW)
}
pt_vm_group_bin_0071 {
0x0: frame_vm_group_bin_2875 (RW)
0x100: frame_vm_group_bin_8865 (RW)
0x101: frame_vm_group_bin_1677 (RW)
0x102: frame_vm_group_bin_17794 (RW)
0x103: frame_vm_group_bin_10685 (RW)
0x104: frame_vm_group_bin_3503 (RW)
0x105: frame_vm_group_bin_19608 (RW)
0x106: frame_vm_group_bin_12428 (RW)
0x107: frame_vm_group_bin_5338 (RW)
0x108: frame_vm_group_bin_21433 (RW)
0x109: frame_vm_group_bin_14257 (RW)
0x10: frame_vm_group_bin_4710 (RW)
0x10a: frame_vm_group_bin_7044 (RW)
0x10b: frame_vm_group_bin_23248 (RW)
0x10c: frame_vm_group_bin_16091 (RW)
0x10d: frame_vm_group_bin_8897 (RW)
0x10e: frame_vm_group_bin_1709 (RW)
0x10f: frame_vm_group_bin_17824 (RW)
0x110: frame_vm_group_bin_10717 (RW)
0x111: frame_vm_group_bin_3531 (RW)
0x112: frame_vm_group_bin_19639 (RW)
0x113: frame_vm_group_bin_12459 (RW)
0x114: frame_vm_group_bin_5369 (RW)
0x115: frame_vm_group_bin_21465 (RW)
0x116: frame_vm_group_bin_14289 (RW)
0x117: frame_vm_group_bin_7075 (RW)
0x118: frame_vm_group_bin_17913 (RW)
0x119: frame_vm_group_bin_16123 (RW)
0x11: frame_vm_group_bin_20832 (RW)
0x11a: frame_vm_group_bin_8930 (RW)
0x11b: frame_vm_group_bin_1742 (RW)
0x11c: frame_vm_group_bin_17853 (RW)
0x11d: frame_vm_group_bin_10750 (RW)
0x11e: frame_vm_group_bin_3563 (RW)
0x11f: frame_vm_group_bin_19667 (RW)
0x120: frame_vm_group_bin_12492 (RW)
0x121: frame_vm_group_bin_5402 (RW)
0x122: frame_vm_group_bin_21497 (RW)
0x123: frame_vm_group_bin_14321 (RW)
0x124: frame_vm_group_bin_7107 (RW)
0x125: frame_vm_group_bin_22647 (RW)
0x126: frame_vm_group_bin_16155 (RW)
0x127: frame_vm_group_bin_8962 (RW)
0x128: frame_vm_group_bin_1774 (RW)
0x129: frame_vm_group_bin_17878 (RW)
0x12: frame_vm_group_bin_13634 (RW)
0x12a: frame_vm_group_bin_10782 (RW)
0x12b: frame_vm_group_bin_3597 (RW)
0x12c: frame_vm_group_bin_19697 (RW)
0x12d: frame_vm_group_bin_12525 (RW)
0x12e: frame_vm_group_bin_5435 (RW)
0x12f: frame_vm_group_bin_21530 (RW)
0x130: frame_vm_group_bin_14354 (RW)
0x131: frame_vm_group_bin_7139 (RW)
0x132: frame_vm_group_bin_0058 (RW)
0x133: frame_vm_group_bin_16188 (RW)
0x134: frame_vm_group_bin_8995 (RW)
0x135: frame_vm_group_bin_1807 (RW)
0x136: frame_vm_group_bin_21562 (RW)
0x137: frame_vm_group_bin_10815 (RW)
0x138: frame_vm_group_bin_3630 (RW)
0x139: frame_vm_group_bin_19730 (RW)
0x13: frame_vm_group_bin_6444 (RW)
0x13a: frame_vm_group_bin_12559 (RW)
0x13b: frame_vm_group_bin_5468 (RW)
0x13c: frame_vm_group_bin_21564 (RW)
0x13d: frame_vm_group_bin_14388 (RW)
0x13e: frame_vm_group_bin_7175 (RW)
0x13f: frame_vm_group_bin_8646 (RW)
0x140: frame_vm_group_bin_16219 (RW)
0x141: frame_vm_group_bin_9029 (RW)
0x142: frame_vm_group_bin_1841 (RW)
0x143: frame_vm_group_bin_17942 (RW)
0x144: frame_vm_group_bin_10849 (RW)
0x145: frame_vm_group_bin_3664 (RW)
0x146: frame_vm_group_bin_19764 (RW)
0x147: frame_vm_group_bin_12592 (RW)
0x148: frame_vm_group_bin_5500 (RW)
0x149: frame_vm_group_bin_21597 (RW)
0x14: frame_vm_group_bin_22641 (RW)
0x14a: frame_vm_group_bin_14421 (RW)
0x14b: frame_vm_group_bin_7208 (RW)
0x14c: frame_vm_group_bin_0110 (RW)
0x14d: frame_vm_group_bin_16245 (RW)
0x14e: frame_vm_group_bin_9062 (RW)
0x14f: frame_vm_group_bin_1874 (RW)
0x150: frame_vm_group_bin_7549 (RW)
0x151: frame_vm_group_bin_10881 (RW)
0x152: frame_vm_group_bin_3697 (RW)
0x153: frame_vm_group_bin_19797 (RW)
0x154: frame_vm_group_bin_12625 (RW)
0x155: frame_vm_group_bin_5532 (RW)
0x156: frame_vm_group_bin_21630 (RW)
0x157: frame_vm_group_bin_14454 (RW)
0x158: frame_vm_group_bin_7241 (RW)
0x159: frame_vm_group_bin_0132 (RW)
0x15: frame_vm_group_bin_15459 (RW)
0x15a: frame_vm_group_bin_16273 (RW)
0x15b: frame_vm_group_bin_9096 (RW)
0x15c: frame_vm_group_bin_1908 (RW)
0x15d: frame_vm_group_bin_18006 (RW)
0x15e: frame_vm_group_bin_10916 (RW)
0x15f: frame_vm_group_bin_3731 (RW)
0x160: frame_vm_group_bin_19831 (RW)
0x161: frame_vm_group_bin_12657 (RW)
0x162: frame_vm_group_bin_5566 (RW)
0x163: frame_vm_group_bin_21664 (RW)
0x164: frame_vm_group_bin_14488 (RW)
0x165: frame_vm_group_bin_7275 (RW)
0x166: frame_vm_group_bin_22670 (RW)
0x167: frame_vm_group_bin_16304 (RW)
0x168: frame_vm_group_bin_9129 (RW)
0x169: frame_vm_group_bin_1941 (RW)
0x16: frame_vm_group_bin_8268 (RW)
0x16a: frame_vm_group_bin_18039 (RW)
0x16b: frame_vm_group_bin_10949 (RW)
0x16c: frame_vm_group_bin_3764 (RW)
0x16d: frame_vm_group_bin_19864 (RW)
0x16e: frame_vm_group_bin_12681 (RW)
0x16f: frame_vm_group_bin_5598 (RW)
0x170: frame_vm_group_bin_21696 (RW)
0x171: frame_vm_group_bin_14522 (RW)
0x172: frame_vm_group_bin_7307 (RW)
0x173: frame_vm_group_bin_0182 (RW)
0x174: frame_vm_group_bin_16336 (RW)
0x175: frame_vm_group_bin_9161 (RW)
0x176: frame_vm_group_bin_1973 (RW)
0x177: frame_vm_group_bin_18071 (RW)
0x178: frame_vm_group_bin_10981 (RW)
0x179: frame_vm_group_bin_3796 (RW)
0x17: frame_vm_group_bin_1083 (RW)
0x17a: frame_vm_group_bin_19897 (RW)
0x17b: frame_vm_group_bin_12706 (RW)
0x17c: frame_vm_group_bin_5630 (RW)
0x17d: frame_vm_group_bin_21730 (RW)
0x17e: frame_vm_group_bin_14556 (RW)
0x17f: frame_vm_group_bin_7341 (RW)
0x180: frame_vm_group_bin_0214 (RW)
0x181: frame_vm_group_bin_16370 (RW)
0x182: frame_vm_group_bin_9193 (RW)
0x183: frame_vm_group_bin_2007 (RW)
0x184: frame_vm_group_bin_18103 (RW)
0x185: frame_vm_group_bin_11015 (RW)
0x186: frame_vm_group_bin_3830 (RW)
0x187: frame_vm_group_bin_19928 (RW)
0x188: frame_vm_group_bin_12732 (RW)
0x189: frame_vm_group_bin_5663 (RW)
0x18: frame_vm_group_bin_17304 (RW)
0x18a: frame_vm_group_bin_21763 (RW)
0x18b: frame_vm_group_bin_14589 (RW)
0x18c: frame_vm_group_bin_7374 (RW)
0x18d: frame_vm_group_bin_13310 (RW)
0x18e: frame_vm_group_bin_16403 (RW)
0x18f: frame_vm_group_bin_9220 (RW)
0x190: frame_vm_group_bin_2040 (RW)
0x191: frame_vm_group_bin_18136 (RW)
0x192: frame_vm_group_bin_11048 (RW)
0x193: frame_vm_group_bin_3863 (RW)
0x194: frame_vm_group_bin_19961 (RW)
0x195: frame_vm_group_bin_12760 (RW)
0x196: frame_vm_group_bin_5696 (RW)
0x197: frame_vm_group_bin_21795 (RW)
0x198: frame_vm_group_bin_14621 (RW)
0x199: frame_vm_group_bin_7407 (RW)
0x19: frame_vm_group_bin_10098 (RW)
0x19a: frame_vm_group_bin_17958 (RW)
0x19b: frame_vm_group_bin_16437 (RW)
0x19c: frame_vm_group_bin_9245 (RW)
0x19d: frame_vm_group_bin_2074 (RW)
0x19e: frame_vm_group_bin_18170 (RW)
0x19f: frame_vm_group_bin_11082 (RW)
0x1: frame_vm_group_bin_18947 (RW)
0x1a0: frame_vm_group_bin_3897 (RW)
0x1a1: frame_vm_group_bin_19993 (RW)
0x1a2: frame_vm_group_bin_12794 (RW)
0x1a3: frame_vm_group_bin_5730 (RW)
0x1a4: frame_vm_group_bin_21830 (RW)
0x1a5: frame_vm_group_bin_14655 (RW)
0x1a6: frame_vm_group_bin_7441 (RW)
0x1a7: frame_vm_group_bin_22693 (RW)
0x1a8: frame_vm_group_bin_16470 (RW)
0x1a9: frame_vm_group_bin_9268 (RW)
0x1a: frame_vm_group_bin_2942 (RW)
0x1aa: frame_vm_group_bin_2107 (RW)
0x1ab: frame_vm_group_bin_18202 (RW)
0x1ac: frame_vm_group_bin_11115 (RW)
0x1ad: frame_vm_group_bin_3930 (RW)
0x1ae: frame_vm_group_bin_20026 (RW)
0x1af: frame_vm_group_bin_12826 (RW)
0x1b0: frame_vm_group_bin_5756 (RW)
0x1b1: frame_vm_group_bin_21863 (RW)
0x1b2: frame_vm_group_bin_14688 (RW)
0x1b3: frame_vm_group_bin_7474 (RW)
0x1b4: frame_vm_group_bin_0321 (RW)
0x1b5: frame_vm_group_bin_16503 (RW)
0x1b6: frame_vm_group_bin_9294 (RW)
0x1b7: frame_vm_group_bin_2141 (RW)
0x1b8: frame_vm_group_bin_18235 (RW)
0x1b9: frame_vm_group_bin_11147 (RW)
0x1b: frame_vm_group_bin_19012 (RW)
0x1ba: frame_vm_group_bin_3963 (RW)
0x1bb: frame_vm_group_bin_20060 (RW)
0x1bc: frame_vm_group_bin_12860 (RW)
0x1bd: frame_vm_group_bin_5781 (RW)
0x1be: frame_vm_group_bin_21897 (RW)
0x1bf: frame_vm_group_bin_14722 (RW)
0x1c0: frame_vm_group_bin_7507 (RW)
0x1c1: frame_vm_group_bin_0353 (RW)
0x1c2: frame_vm_group_bin_16537 (RW)
0x1c3: frame_vm_group_bin_9325 (RW)
0x1c4: frame_vm_group_bin_2175 (RW)
0x1c5: frame_vm_group_bin_18269 (RW)
0x1c6: frame_vm_group_bin_11181 (RW)
0x1c7: frame_vm_group_bin_3996 (RW)
0x1c8: frame_vm_group_bin_20093 (RW)
0x1c9: frame_vm_group_bin_12893 (RW)
0x1c: frame_vm_group_bin_11866 (RW)
0x1ca: frame_vm_group_bin_7170 (RW)
0x1cb: frame_vm_group_bin_21929 (RW)
0x1cc: frame_vm_group_bin_14754 (RW)
0x1cd: frame_vm_group_bin_7539 (RW)
0x1ce: frame_vm_group_bin_13334 (RW)
0x1cf: frame_vm_group_bin_16569 (RW)
0x1d0: frame_vm_group_bin_9358 (RW)
0x1d1: frame_vm_group_bin_2206 (RW)
0x1d2: frame_vm_group_bin_18302 (RW)
0x1d3: frame_vm_group_bin_11214 (RW)
0x1d4: frame_vm_group_bin_4029 (RW)
0x1d5: frame_vm_group_bin_20125 (RW)
0x1d6: frame_vm_group_bin_12926 (RW)
0x1d7: frame_vm_group_bin_0435 (RW)
0x1d8: frame_vm_group_bin_21962 (RW)
0x1d9: frame_vm_group_bin_14786 (RW)
0x1d: frame_vm_group_bin_4743 (RW)
0x1da: frame_vm_group_bin_7572 (RW)
0x1db: frame_vm_group_bin_0414 (RW)
0x1dc: frame_vm_group_bin_16602 (RW)
0x1dd: frame_vm_group_bin_9393 (RW)
0x1de: frame_vm_group_bin_2235 (RW)
0x1df: frame_vm_group_bin_18336 (RW)
0x1e0: frame_vm_group_bin_11248 (RW)
0x1e1: frame_vm_group_bin_4063 (RW)
0x1e2: frame_vm_group_bin_20158 (RW)
0x1e3: frame_vm_group_bin_12959 (RW)
0x1e4: frame_vm_group_bin_5163 (RW)
0x1e5: frame_vm_group_bin_21996 (RW)
0x1e6: frame_vm_group_bin_14820 (RW)
0x1e7: frame_vm_group_bin_7605 (RW)
0x1e8: frame_vm_group_bin_0445 (RW)
0x1e9: frame_vm_group_bin_16635 (RW)
0x1e: frame_vm_group_bin_20861 (RW)
0x1ea: frame_vm_group_bin_9426 (RW)
0x1eb: frame_vm_group_bin_2266 (RW)
0x1ec: frame_vm_group_bin_18369 (RW)
0x1ed: frame_vm_group_bin_11281 (RW)
0x1ee: frame_vm_group_bin_4096 (RW)
0x1ef: frame_vm_group_bin_20190 (RW)
0x1f0: frame_vm_group_bin_12992 (RW)
0x1f1: frame_vm_group_bin_9793 (RW)
0x1f2: frame_vm_group_bin_22025 (RW)
0x1f3: frame_vm_group_bin_14853 (RW)
0x1f4: frame_vm_group_bin_7638 (RW)
0x1f5: frame_vm_group_bin_0478 (RW)
0x1f6: frame_vm_group_bin_16668 (RW)
0x1f7: frame_vm_group_bin_9459 (RW)
0x1f8: frame_vm_group_bin_2299 (RW)
0x1f9: frame_vm_group_bin_18401 (RW)
0x1f: frame_vm_group_bin_13667 (RW)
0x1fa: frame_vm_group_bin_11315 (RW)
0x1fb: frame_vm_group_bin_4129 (RW)
0x1fc: frame_vm_group_bin_20224 (RW)
0x1fd: frame_vm_group_bin_13028 (RW)
0x1fe: frame_vm_group_bin_5901 (RW)
0x1ff: frame_vm_group_bin_22048 (RW)
0x20: frame_vm_group_bin_6478 (RW)
0x21: frame_vm_group_bin_22675 (RW)
0x22: frame_vm_group_bin_15493 (RW)
0x23: frame_vm_group_bin_8301 (RW)
0x24: frame_vm_group_bin_1113 (RW)
0x25: frame_vm_group_bin_17338 (RW)
0x26: frame_vm_group_bin_10132 (RW)
0x27: frame_vm_group_bin_2975 (RW)
0x28: frame_vm_group_bin_19045 (RW)
0x29: frame_vm_group_bin_11103 (RW)
0x2: frame_vm_group_bin_11804 (RW)
0x2a: frame_vm_group_bin_4776 (RW)
0x2b: frame_vm_group_bin_20885 (RW)
0x2c: frame_vm_group_bin_13700 (RW)
0x2d: frame_vm_group_bin_6511 (RW)
0x2e: frame_vm_group_bin_22708 (RW)
0x2f: frame_vm_group_bin_15525 (RW)
0x30: frame_vm_group_bin_8334 (RW)
0x31: frame_vm_group_bin_1145 (RW)
0x32: frame_vm_group_bin_17370 (RW)
0x33: frame_vm_group_bin_10167 (RW)
0x34: frame_vm_group_bin_3008 (RW)
0x35: frame_vm_group_bin_19078 (RW)
0x36: frame_vm_group_bin_11917 (RW)
0x37: frame_vm_group_bin_4809 (RW)
0x38: frame_vm_group_bin_20913 (RW)
0x39: frame_vm_group_bin_13732 (RW)
0x3: frame_vm_group_bin_4678 (RW)
0x3a: frame_vm_group_bin_6545 (RW)
0x3b: frame_vm_group_bin_22742 (RW)
0x3c: frame_vm_group_bin_15558 (RW)
0x3d: frame_vm_group_bin_8368 (RW)
0x3e: frame_vm_group_bin_1179 (RW)
0x3f: frame_vm_group_bin_17401 (RW)
0x40: frame_vm_group_bin_10201 (RW)
0x41: frame_vm_group_bin_3042 (RW)
0x42: frame_vm_group_bin_19111 (RW)
0x43: frame_vm_group_bin_11947 (RW)
0x44: frame_vm_group_bin_4842 (RW)
0x45: frame_vm_group_bin_20943 (RW)
0x46: frame_vm_group_bin_13767 (RW)
0x47: frame_vm_group_bin_6578 (RW)
0x48: frame_vm_group_bin_22774 (RW)
0x49: frame_vm_group_bin_15591 (RW)
0x4: frame_vm_group_bin_20800 (RW)
0x4a: frame_vm_group_bin_8401 (RW)
0x4b: frame_vm_group_bin_1212 (RW)
0x4c: frame_vm_group_bin_17426 (RW)
0x4d: frame_vm_group_bin_10234 (RW)
0x4e: frame_vm_group_bin_3075 (RW)
0x4f: frame_vm_group_bin_19143 (RW)
0x50: frame_vm_group_bin_11980 (RW)
0x51: frame_vm_group_bin_4875 (RW)
0x52: frame_vm_group_bin_20968 (RW)
0x53: frame_vm_group_bin_13800 (RW)
0x54: frame_vm_group_bin_6611 (RW)
0x55: frame_vm_group_bin_22807 (RW)
0x56: frame_vm_group_bin_15624 (RW)
0x57: frame_vm_group_bin_8434 (RW)
0x58: frame_vm_group_bin_1245 (RW)
0x59: frame_vm_group_bin_18095 (RW)
0x5: frame_vm_group_bin_13601 (RW)
0x5a: frame_vm_group_bin_10268 (RW)
0x5b: frame_vm_group_bin_3109 (RW)
0x5c: frame_vm_group_bin_19177 (RW)
0x5d: frame_vm_group_bin_12013 (RW)
0x5e: frame_vm_group_bin_4909 (RW)
0x5f: frame_vm_group_bin_21002 (RW)
0x60: frame_vm_group_bin_13832 (RW)
0x61: frame_vm_group_bin_6645 (RW)
0x62: frame_vm_group_bin_22841 (RW)
0x63: frame_vm_group_bin_15658 (RW)
0x64: frame_vm_group_bin_8468 (RW)
0x65: frame_vm_group_bin_1276 (RW)
0x66: frame_vm_group_bin_2869 (RW)
0x67: frame_vm_group_bin_10301 (RW)
0x68: frame_vm_group_bin_3141 (RW)
0x69: frame_vm_group_bin_19210 (RW)
0x6: frame_vm_group_bin_6411 (RW)
0x6a: frame_vm_group_bin_11125 (RW)
0x6b: frame_vm_group_bin_4940 (RW)
0x6c: frame_vm_group_bin_21035 (RW)
0x6d: frame_vm_group_bin_13861 (RW)
0x6e: frame_vm_group_bin_6678 (RW)
0x6f: frame_vm_group_bin_22874 (RW)
0x70: frame_vm_group_bin_15691 (RW)
0x71: frame_vm_group_bin_8501 (RW)
0x72: frame_vm_group_bin_1309 (RW)
0x73: frame_vm_group_bin_21492 (RW)
0x74: frame_vm_group_bin_10334 (RW)
0x75: frame_vm_group_bin_3174 (RW)
0x76: frame_vm_group_bin_19243 (RW)
0x77: frame_vm_group_bin_12070 (RW)
0x78: frame_vm_group_bin_4971 (RW)
0x79: frame_vm_group_bin_21069 (RW)
0x7: frame_vm_group_bin_22608 (RW)
0x7a: frame_vm_group_bin_13892 (RW)
0x7b: frame_vm_group_bin_6712 (RW)
0x7c: frame_vm_group_bin_22908 (RW)
0x7d: frame_vm_group_bin_15725 (RW)
0x7e: frame_vm_group_bin_8534 (RW)
0x7f: frame_vm_group_bin_1342 (RW)
0x80: frame_vm_group_bin_2871 (RW)
0x81: frame_vm_group_bin_10368 (RW)
0x82: frame_vm_group_bin_3208 (RW)
0x83: frame_vm_group_bin_19277 (RW)
0x84: frame_vm_group_bin_12104 (RW)
0x85: frame_vm_group_bin_5005 (RW)
0x86: frame_vm_group_bin_21103 (RW)
0x87: frame_vm_group_bin_13925 (RW)
0x88: frame_vm_group_bin_6744 (RW)
0x89: frame_vm_group_bin_22941 (RW)
0x8: frame_vm_group_bin_15426 (RW)
0x8a: frame_vm_group_bin_15758 (RW)
0x8b: frame_vm_group_bin_8565 (RW)
0x8c: frame_vm_group_bin_1376 (RW)
0x8d: frame_vm_group_bin_7481 (RW)
0x8e: frame_vm_group_bin_10397 (RW)
0x8f: frame_vm_group_bin_3240 (RW)
0x90: frame_vm_group_bin_19310 (RW)
0x91: frame_vm_group_bin_12136 (RW)
0x92: frame_vm_group_bin_5038 (RW)
0x93: frame_vm_group_bin_21136 (RW)
0x94: frame_vm_group_bin_13958 (RW)
0x95: frame_vm_group_bin_6776 (RW)
0x96: frame_vm_group_bin_22973 (RW)
0x97: frame_vm_group_bin_15791 (RW)
0x98: frame_vm_group_bin_8598 (RW)
0x99: frame_vm_group_bin_1409 (RW)
0x9: frame_vm_group_bin_8235 (RW)
0x9a: frame_vm_group_bin_12143 (RW)
0x9b: frame_vm_group_bin_10424 (RW)
0x9c: frame_vm_group_bin_3274 (RW)
0x9d: frame_vm_group_bin_19344 (RW)
0x9e: frame_vm_group_bin_12167 (RW)
0x9f: frame_vm_group_bin_5073 (RW)
0xa0: frame_vm_group_bin_21169 (RW)
0xa1: frame_vm_group_bin_13992 (RW)
0xa2: frame_vm_group_bin_6809 (RW)
0xa3: frame_vm_group_bin_23006 (RW)
0xa4: frame_vm_group_bin_15823 (RW)
0xa5: frame_vm_group_bin_8631 (RW)
0xa6: frame_vm_group_bin_1443 (RW)
0xa7: frame_vm_group_bin_16884 (RW)
0xa8: frame_vm_group_bin_10454 (RW)
0xa9: frame_vm_group_bin_3307 (RW)
0xa: frame_vm_group_bin_1059 (RW)
0xaa: frame_vm_group_bin_19377 (RW)
0xab: frame_vm_group_bin_12199 (RW)
0xac: frame_vm_group_bin_5106 (RW)
0xad: frame_vm_group_bin_21202 (RW)
0xae: frame_vm_group_bin_14025 (RW)
0xaf: frame_vm_group_bin_6838 (RW)
0xb0: frame_vm_group_bin_23039 (RW)
0xb1: frame_vm_group_bin_15856 (RW)
0xb2: frame_vm_group_bin_8664 (RW)
0xb3: frame_vm_group_bin_1476 (RW)
0xb4: frame_vm_group_bin_17616 (RW)
0xb5: frame_vm_group_bin_10487 (RW)
0xb6: frame_vm_group_bin_3340 (RW)
0xb7: frame_vm_group_bin_19410 (RW)
0xb8: frame_vm_group_bin_12229 (RW)
0xb9: frame_vm_group_bin_5139 (RW)
0xb: frame_vm_group_bin_17271 (RW)
0xba: frame_vm_group_bin_21236 (RW)
0xbb: frame_vm_group_bin_14059 (RW)
0xbc: frame_vm_group_bin_6866 (RW)
0xbd: frame_vm_group_bin_23073 (RW)
0xbe: frame_vm_group_bin_15890 (RW)
0xbf: frame_vm_group_bin_8699 (RW)
0xc0: frame_vm_group_bin_1510 (RW)
0xc1: frame_vm_group_bin_17650 (RW)
0xc2: frame_vm_group_bin_10520 (RW)
0xc3: frame_vm_group_bin_0045 (RW)
0xc4: frame_vm_group_bin_19441 (RW)
0xc5: frame_vm_group_bin_12262 (RW)
0xc6: frame_vm_group_bin_5173 (RW)
0xc7: frame_vm_group_bin_21269 (RW)
0xc8: frame_vm_group_bin_14092 (RW)
0xc9: frame_vm_group_bin_6891 (RW)
0xc: frame_vm_group_bin_10065 (RW)
0xca: frame_vm_group_bin_23106 (RW)
0xcb: frame_vm_group_bin_15923 (RW)
0xcc: frame_vm_group_bin_8732 (RW)
0xcd: frame_vm_group_bin_1543 (RW)
0xce: frame_vm_group_bin_7504 (RW)
0xcf: frame_vm_group_bin_10553 (RW)
0xd0: frame_vm_group_bin_3402 (RW)
0xd1: frame_vm_group_bin_19473 (RW)
0xd2: frame_vm_group_bin_12295 (RW)
0xd3: frame_vm_group_bin_5206 (RW)
0xd4: frame_vm_group_bin_21302 (RW)
0xd5: frame_vm_group_bin_14125 (RW)
0xd6: frame_vm_group_bin_6915 (RW)
0xd7: frame_vm_group_bin_23139 (RW)
0xd8: frame_vm_group_bin_15956 (RW)
0xd9: frame_vm_group_bin_8765 (RW)
0xd: frame_vm_group_bin_2908 (RW)
0xda: frame_vm_group_bin_1577 (RW)
0xdb: frame_vm_group_bin_17710 (RW)
0xdc: frame_vm_group_bin_10587 (RW)
0xdd: frame_vm_group_bin_3427 (RW)
0xde: frame_vm_group_bin_19507 (RW)
0xdf: frame_vm_group_bin_12328 (RW)
0xe0: frame_vm_group_bin_5240 (RW)
0xe1: frame_vm_group_bin_21334 (RW)
0xe2: frame_vm_group_bin_14159 (RW)
0xe3: frame_vm_group_bin_6946 (RW)
0xe4: frame_vm_group_bin_23172 (RW)
0xe5: frame_vm_group_bin_15992 (RW)
0xe6: frame_vm_group_bin_8799 (RW)
0xe7: frame_vm_group_bin_1610 (RW)
0xe8: frame_vm_group_bin_17736 (RW)
0xe9: frame_vm_group_bin_10620 (RW)
0xe: frame_vm_group_bin_18978 (RW)
0xea: frame_vm_group_bin_3449 (RW)
0xeb: frame_vm_group_bin_19540 (RW)
0xec: frame_vm_group_bin_12361 (RW)
0xed: frame_vm_group_bin_5273 (RW)
0xee: frame_vm_group_bin_21367 (RW)
0xef: frame_vm_group_bin_14191 (RW)
0xf0: frame_vm_group_bin_6978 (RW)
0xf1: frame_vm_group_bin_23203 (RW)
0xf2: frame_vm_group_bin_16025 (RW)
0xf3: frame_vm_group_bin_8832 (RW)
0xf4: frame_vm_group_bin_1643 (RW)
0xf5: frame_vm_group_bin_17763 (RW)
0xf6: frame_vm_group_bin_10652 (RW)
0xf7: frame_vm_group_bin_3475 (RW)
0xf8: frame_vm_group_bin_19573 (RW)
0xf9: frame_vm_group_bin_12394 (RW)
0xf: frame_vm_group_bin_11836 (RW)
0xfa: frame_vm_group_bin_5307 (RW)
0xfb: frame_vm_group_bin_21401 (RW)
0xfc: frame_vm_group_bin_14225 (RW)
0xfd: frame_vm_group_bin_7012 (RW)
0xfe: frame_vm_group_bin_23227 (RW)
0xff: frame_vm_group_bin_16059 (RW)
}
pt_vm_group_bin_0079 {
0x0: frame_vm_group_bin_3589 (RW)
0x100: frame_vm_group_bin_9585 (RW)
0x101: frame_vm_group_bin_2424 (RW)
0x102: frame_vm_group_bin_18515 (RW)
0x103: frame_vm_group_bin_11436 (RW)
0x104: frame_vm_group_bin_4252 (RW)
0x105: frame_vm_group_bin_20350 (RW)
0x106: frame_vm_group_bin_13153 (RW)
0x107: frame_vm_group_bin_5998 (RW)
0x108: frame_vm_group_bin_22161 (RW)
0x109: frame_vm_group_bin_15012 (RW)
0x10: frame_vm_group_bin_5459 (RW)
0x10a: frame_vm_group_bin_7796 (RW)
0x10b: frame_vm_group_bin_0630 (RW)
0x10c: frame_vm_group_bin_16827 (RW)
0x10d: frame_vm_group_bin_9618 (RW)
0x10e: frame_vm_group_bin_2457 (RW)
0x10f: frame_vm_group_bin_18540 (RW)
0x110: frame_vm_group_bin_11469 (RW)
0x111: frame_vm_group_bin_4285 (RW)
0x112: frame_vm_group_bin_20383 (RW)
0x113: frame_vm_group_bin_13186 (RW)
0x114: frame_vm_group_bin_6029 (RW)
0x115: frame_vm_group_bin_22194 (RW)
0x116: frame_vm_group_bin_15040 (RW)
0x117: frame_vm_group_bin_7829 (RW)
0x118: frame_vm_group_bin_0664 (RW)
0x119: frame_vm_group_bin_16860 (RW)
0x11: frame_vm_group_bin_21555 (RW)
0x11a: frame_vm_group_bin_9652 (RW)
0x11b: frame_vm_group_bin_2490 (RW)
0x11c: frame_vm_group_bin_18567 (RW)
0x11d: frame_vm_group_bin_11503 (RW)
0x11e: frame_vm_group_bin_4319 (RW)
0x11f: frame_vm_group_bin_20417 (RW)
0x120: frame_vm_group_bin_13220 (RW)
0x121: frame_vm_group_bin_6055 (RW)
0x122: frame_vm_group_bin_22228 (RW)
0x123: frame_vm_group_bin_15068 (RW)
0x124: frame_vm_group_bin_7862 (RW)
0x125: frame_vm_group_bin_0698 (RW)
0x126: frame_vm_group_bin_16892 (RW)
0x127: frame_vm_group_bin_9684 (RW)
0x128: frame_vm_group_bin_2523 (RW)
0x129: frame_vm_group_bin_18600 (RW)
0x12: frame_vm_group_bin_14379 (RW)
0x12a: frame_vm_group_bin_11536 (RW)
0x12b: frame_vm_group_bin_4354 (RW)
0x12c: frame_vm_group_bin_20450 (RW)
0x12d: frame_vm_group_bin_13253 (RW)
0x12e: frame_vm_group_bin_6081 (RW)
0x12f: frame_vm_group_bin_22261 (RW)
0x130: frame_vm_group_bin_15092 (RW)
0x131: frame_vm_group_bin_7895 (RW)
0x132: frame_vm_group_bin_0731 (RW)
0x133: frame_vm_group_bin_16925 (RW)
0x134: frame_vm_group_bin_9717 (RW)
0x135: frame_vm_group_bin_2556 (RW)
0x136: frame_vm_group_bin_18633 (RW)
0x137: frame_vm_group_bin_11566 (RW)
0x138: frame_vm_group_bin_4387 (RW)
0x139: frame_vm_group_bin_20483 (RW)
0x13: frame_vm_group_bin_7164 (RW)
0x13a: frame_vm_group_bin_13287 (RW)
0x13b: frame_vm_group_bin_14386 (RW)
0x13c: frame_vm_group_bin_22294 (RW)
0x13d: frame_vm_group_bin_15120 (RW)
0x13e: frame_vm_group_bin_7930 (RW)
0x13f: frame_vm_group_bin_0765 (RW)
0x140: frame_vm_group_bin_16959 (RW)
0x141: frame_vm_group_bin_9751 (RW)
0x142: frame_vm_group_bin_2590 (RW)
0x143: frame_vm_group_bin_18666 (RW)
0x144: frame_vm_group_bin_11595 (RW)
0x145: frame_vm_group_bin_4421 (RW)
0x146: frame_vm_group_bin_20517 (RW)
0x147: frame_vm_group_bin_13319 (RW)
0x148: frame_vm_group_bin_6144 (RW)
0x149: frame_vm_group_bin_22327 (RW)
0x14: frame_vm_group_bin_0077 (RW)
0x14a: frame_vm_group_bin_15143 (RW)
0x14b: frame_vm_group_bin_7963 (RW)
0x14c: frame_vm_group_bin_0798 (RW)
0x14d: frame_vm_group_bin_16992 (RW)
0x14e: frame_vm_group_bin_9784 (RW)
0x14f: frame_vm_group_bin_2623 (RW)
0x150: frame_vm_group_bin_18699 (RW)
0x151: frame_vm_group_bin_11620 (RW)
0x152: frame_vm_group_bin_4454 (RW)
0x153: frame_vm_group_bin_20550 (RW)
0x154: frame_vm_group_bin_13352 (RW)
0x155: frame_vm_group_bin_6177 (RW)
0x156: frame_vm_group_bin_22359 (RW)
0x157: frame_vm_group_bin_15175 (RW)
0x158: frame_vm_group_bin_7994 (RW)
0x159: frame_vm_group_bin_0830 (RW)
0x15: frame_vm_group_bin_16210 (RW)
0x15a: frame_vm_group_bin_17026 (RW)
0x15b: frame_vm_group_bin_9818 (RW)
0x15c: frame_vm_group_bin_2657 (RW)
0x15d: frame_vm_group_bin_18732 (RW)
0x15e: frame_vm_group_bin_10841 (RW)
0x15f: frame_vm_group_bin_4488 (RW)
0x160: frame_vm_group_bin_20584 (RW)
0x161: frame_vm_group_bin_13384 (RW)
0x162: frame_vm_group_bin_5117 (RW)
0x163: frame_vm_group_bin_22393 (RW)
0x164: frame_vm_group_bin_15209 (RW)
0x165: frame_vm_group_bin_8025 (RW)
0x166: frame_vm_group_bin_0864 (RW)
0x167: frame_vm_group_bin_17059 (RW)
0x168: frame_vm_group_bin_9851 (RW)
0x169: frame_vm_group_bin_2690 (RW)
0x16: frame_vm_group_bin_9020 (RW)
0x16a: frame_vm_group_bin_18763 (RW)
0x16b: frame_vm_group_bin_15487 (RW)
0x16c: frame_vm_group_bin_4521 (RW)
0x16d: frame_vm_group_bin_20617 (RW)
0x16e: frame_vm_group_bin_13417 (RW)
0x16f: frame_vm_group_bin_6234 (RW)
0x170: frame_vm_group_bin_22425 (RW)
0x171: frame_vm_group_bin_15243 (RW)
0x172: frame_vm_group_bin_8054 (RW)
0x173: frame_vm_group_bin_0897 (RW)
0x174: frame_vm_group_bin_17092 (RW)
0x175: frame_vm_group_bin_9884 (RW)
0x176: frame_vm_group_bin_2723 (RW)
0x177: frame_vm_group_bin_18796 (RW)
0x178: frame_vm_group_bin_11688 (RW)
0x179: frame_vm_group_bin_4553 (RW)
0x17: frame_vm_group_bin_1832 (RW)
0x17a: frame_vm_group_bin_20651 (RW)
0x17b: frame_vm_group_bin_13451 (RW)
0x17c: frame_vm_group_bin_6266 (RW)
0x17d: frame_vm_group_bin_22459 (RW)
0x17e: frame_vm_group_bin_15277 (RW)
0x17f: frame_vm_group_bin_8086 (RW)
0x180: frame_vm_group_bin_0931 (RW)
0x181: frame_vm_group_bin_17126 (RW)
0x182: frame_vm_group_bin_9917 (RW)
0x183: frame_vm_group_bin_2757 (RW)
0x184: frame_vm_group_bin_18831 (RW)
0x185: frame_vm_group_bin_11717 (RW)
0x186: frame_vm_group_bin_4582 (RW)
0x187: frame_vm_group_bin_20683 (RW)
0x188: frame_vm_group_bin_13484 (RW)
0x189: frame_vm_group_bin_6299 (RW)
0x18: frame_vm_group_bin_17934 (RW)
0x18a: frame_vm_group_bin_22492 (RW)
0x18b: frame_vm_group_bin_15309 (RW)
0x18c: frame_vm_group_bin_8118 (RW)
0x18d: frame_vm_group_bin_0964 (RW)
0x18e: frame_vm_group_bin_17158 (RW)
0x18f: frame_vm_group_bin_9948 (RW)
0x190: frame_vm_group_bin_2790 (RW)
0x191: frame_vm_group_bin_18864 (RW)
0x192: frame_vm_group_bin_6135 (RW)
0x193: frame_vm_group_bin_4604 (RW)
0x194: frame_vm_group_bin_20716 (RW)
0x195: frame_vm_group_bin_13517 (RW)
0x196: frame_vm_group_bin_6331 (RW)
0x197: frame_vm_group_bin_22525 (RW)
0x198: frame_vm_group_bin_15342 (RW)
0x199: frame_vm_group_bin_8151 (RW)
0x19: frame_vm_group_bin_10840 (RW)
0x19a: frame_vm_group_bin_0998 (RW)
0x19b: frame_vm_group_bin_17191 (RW)
0x19c: frame_vm_group_bin_9982 (RW)
0x19d: frame_vm_group_bin_2824 (RW)
0x19e: frame_vm_group_bin_18898 (RW)
0x19f: frame_vm_group_bin_10865 (RW)
0x1: frame_vm_group_bin_19689 (RW)
0x1a0: frame_vm_group_bin_4630 (RW)
0x1a1: frame_vm_group_bin_20750 (RW)
0x1a2: frame_vm_group_bin_13551 (RW)
0x1a3: frame_vm_group_bin_6365 (RW)
0x1a4: frame_vm_group_bin_22558 (RW)
0x1a5: frame_vm_group_bin_15376 (RW)
0x1a6: frame_vm_group_bin_8185 (RW)
0x1a7: frame_vm_group_bin_1026 (RW)
0x1a8: frame_vm_group_bin_17222 (RW)
0x1a9: frame_vm_group_bin_10015 (RW)
0x1a: frame_vm_group_bin_3656 (RW)
0x1aa: frame_vm_group_bin_2856 (RW)
0x1ab: frame_vm_group_bin_18931 (RW)
0x1ac: frame_vm_group_bin_11788 (RW)
0x1ad: frame_vm_group_bin_4662 (RW)
0x1ae: frame_vm_group_bin_20783 (RW)
0x1af: frame_vm_group_bin_13584 (RW)
0x1b0: frame_vm_group_bin_6395 (RW)
0x1b1: frame_vm_group_bin_22591 (RW)
0x1b2: frame_vm_group_bin_15409 (RW)
0x1b3: frame_vm_group_bin_8218 (RW)
0x1b4: frame_vm_group_bin_1048 (RW)
0x1b5: frame_vm_group_bin_17254 (RW)
0x1b6: frame_vm_group_bin_10048 (RW)
0x1b7: frame_vm_group_bin_2891 (RW)
0x1b8: frame_vm_group_bin_18963 (RW)
0x1b9: frame_vm_group_bin_11820 (RW)
0x1b: frame_vm_group_bin_19756 (RW)
0x1ba: frame_vm_group_bin_4695 (RW)
0x1bb: frame_vm_group_bin_20817 (RW)
0x1bc: frame_vm_group_bin_13618 (RW)
0x1bd: frame_vm_group_bin_6428 (RW)
0x1be: frame_vm_group_bin_22625 (RW)
0x1bf: frame_vm_group_bin_15443 (RW)
0x1c0: frame_vm_group_bin_8252 (RW)
0x1c1: frame_vm_group_bin_1072 (RW)
0x1c2: frame_vm_group_bin_17288 (RW)
0x1c3: frame_vm_group_bin_10082 (RW)
0x1c4: frame_vm_group_bin_2925 (RW)
0x1c5: frame_vm_group_bin_18995 (RW)
0x1c6: frame_vm_group_bin_11851 (RW)
0x1c7: frame_vm_group_bin_4726 (RW)
0x1c8: frame_vm_group_bin_20847 (RW)
0x1c9: frame_vm_group_bin_13650 (RW)
0x1c: frame_vm_group_bin_12584 (RW)
0x1ca: frame_vm_group_bin_6461 (RW)
0x1cb: frame_vm_group_bin_22658 (RW)
0x1cc: frame_vm_group_bin_15476 (RW)
0x1cd: frame_vm_group_bin_8284 (RW)
0x1ce: frame_vm_group_bin_1098 (RW)
0x1cf: frame_vm_group_bin_17321 (RW)
0x1d0: frame_vm_group_bin_10115 (RW)
0x1d1: frame_vm_group_bin_2958 (RW)
0x1d2: frame_vm_group_bin_19028 (RW)
0x1d3: frame_vm_group_bin_6159 (RW)
0x1d4: frame_vm_group_bin_4759 (RW)
0x1d5: frame_vm_group_bin_20871 (RW)
0x1d6: frame_vm_group_bin_13683 (RW)
0x1d7: frame_vm_group_bin_6494 (RW)
0x1d8: frame_vm_group_bin_22691 (RW)
0x1d9: frame_vm_group_bin_15509 (RW)
0x1d: frame_vm_group_bin_5492 (RW)
0x1da: frame_vm_group_bin_8318 (RW)
0x1db: frame_vm_group_bin_1129 (RW)
0x1dc: frame_vm_group_bin_17355 (RW)
0x1dd: frame_vm_group_bin_10151 (RW)
0x1de: frame_vm_group_bin_2992 (RW)
0x1df: frame_vm_group_bin_19062 (RW)
0x1e0: frame_vm_group_bin_10889 (RW)
0x1e1: frame_vm_group_bin_4793 (RW)
0x1e2: frame_vm_group_bin_20901 (RW)
0x1e3: frame_vm_group_bin_13716 (RW)
0x1e4: frame_vm_group_bin_6528 (RW)
0x1e5: frame_vm_group_bin_22725 (RW)
0x1e6: frame_vm_group_bin_15541 (RW)
0x1e7: frame_vm_group_bin_8351 (RW)
0x1e8: frame_vm_group_bin_1162 (RW)
0x1e9: frame_vm_group_bin_17386 (RW)
0x1e: frame_vm_group_bin_21589 (RW)
0x1ea: frame_vm_group_bin_10184 (RW)
0x1eb: frame_vm_group_bin_3025 (RW)
0x1ec: frame_vm_group_bin_19095 (RW)
0x1ed: frame_vm_group_bin_11933 (RW)
0x1ee: frame_vm_group_bin_4825 (RW)
0x1ef: frame_vm_group_bin_20926 (RW)
0x1f0: frame_vm_group_bin_13749 (RW)
0x1f1: frame_vm_group_bin_6561 (RW)
0x1f2: frame_vm_group_bin_22757 (RW)
0x1f3: frame_vm_group_bin_15574 (RW)
0x1f4: frame_vm_group_bin_8384 (RW)
0x1f5: frame_vm_group_bin_1195 (RW)
0x1f6: frame_vm_group_bin_17412 (RW)
0x1f7: frame_vm_group_bin_10217 (RW)
0x1f8: frame_vm_group_bin_3058 (RW)
0x1f9: frame_vm_group_bin_19127 (RW)
0x1f: frame_vm_group_bin_14413 (RW)
0x1fa: frame_vm_group_bin_11964 (RW)
0x1fb: frame_vm_group_bin_4859 (RW)
0x1fc: frame_vm_group_bin_20954 (RW)
0x1fd: frame_vm_group_bin_13784 (RW)
0x1fe: frame_vm_group_bin_6595 (RW)
0x1ff: frame_vm_group_bin_22791 (RW)
0x20: frame_vm_group_bin_7200 (RW)
0x21: frame_vm_group_bin_22551 (RW)
0x22: frame_vm_group_bin_16239 (RW)
0x23: frame_vm_group_bin_9054 (RW)
0x24: frame_vm_group_bin_1866 (RW)
0x25: frame_vm_group_bin_17966 (RW)
0x26: frame_vm_group_bin_10873 (RW)
0x27: frame_vm_group_bin_3689 (RW)
0x28: frame_vm_group_bin_19789 (RW)
0x29: frame_vm_group_bin_12617 (RW)
0x2: frame_vm_group_bin_12517 (RW)
0x2a: frame_vm_group_bin_5524 (RW)
0x2b: frame_vm_group_bin_21622 (RW)
0x2c: frame_vm_group_bin_14446 (RW)
0x2d: frame_vm_group_bin_7233 (RW)
0x2e: frame_vm_group_bin_3917 (RW)
0x2f: frame_vm_group_bin_16265 (RW)
0x30: frame_vm_group_bin_9087 (RW)
0x31: frame_vm_group_bin_1899 (RW)
0x32: frame_vm_group_bin_17997 (RW)
0x33: frame_vm_group_bin_10907 (RW)
0x34: frame_vm_group_bin_3722 (RW)
0x35: frame_vm_group_bin_19822 (RW)
0x36: frame_vm_group_bin_12648 (RW)
0x37: frame_vm_group_bin_5557 (RW)
0x38: frame_vm_group_bin_21655 (RW)
0x39: frame_vm_group_bin_14479 (RW)
0x3: frame_vm_group_bin_5427 (RW)
0x3a: frame_vm_group_bin_7267 (RW)
0x3b: frame_vm_group_bin_8554 (RW)
0x3c: frame_vm_group_bin_16296 (RW)
0x3d: frame_vm_group_bin_9121 (RW)
0x3e: frame_vm_group_bin_1933 (RW)
0x3f: frame_vm_group_bin_18031 (RW)
0x40: frame_vm_group_bin_10941 (RW)
0x41: frame_vm_group_bin_3756 (RW)
0x42: frame_vm_group_bin_19856 (RW)
0x43: frame_vm_group_bin_12676 (RW)
0x44: frame_vm_group_bin_5590 (RW)
0x45: frame_vm_group_bin_21688 (RW)
0x46: frame_vm_group_bin_14514 (RW)
0x47: frame_vm_group_bin_7299 (RW)
0x48: frame_vm_group_bin_0174 (RW)
0x49: frame_vm_group_bin_16328 (RW)
0x4: frame_vm_group_bin_21522 (RW)
0x4a: frame_vm_group_bin_9153 (RW)
0x4b: frame_vm_group_bin_1965 (RW)
0x4c: frame_vm_group_bin_18063 (RW)
0x4d: frame_vm_group_bin_10973 (RW)
0x4e: frame_vm_group_bin_3788 (RW)
0x4f: frame_vm_group_bin_19888 (RW)
0x50: frame_vm_group_bin_12699 (RW)
0x51: frame_vm_group_bin_5621 (RW)
0x52: frame_vm_group_bin_21721 (RW)
0x53: frame_vm_group_bin_14547 (RW)
0x54: frame_vm_group_bin_7332 (RW)
0x55: frame_vm_group_bin_0206 (RW)
0x56: frame_vm_group_bin_16361 (RW)
0x57: frame_vm_group_bin_9184 (RW)
0x58: frame_vm_group_bin_1998 (RW)
0x59: frame_vm_group_bin_18096 (RW)
0x5: frame_vm_group_bin_14346 (RW)
0x5a: frame_vm_group_bin_11007 (RW)
0x5b: frame_vm_group_bin_3822 (RW)
0x5c: frame_vm_group_bin_19921 (RW)
0x5d: frame_vm_group_bin_12725 (RW)
0x5e: frame_vm_group_bin_5655 (RW)
0x5f: frame_vm_group_bin_21755 (RW)
0x60: frame_vm_group_bin_14581 (RW)
0x61: frame_vm_group_bin_7366 (RW)
0x62: frame_vm_group_bin_22574 (RW)
0x63: frame_vm_group_bin_16395 (RW)
0x64: frame_vm_group_bin_9214 (RW)
0x65: frame_vm_group_bin_2032 (RW)
0x66: frame_vm_group_bin_18128 (RW)
0x67: frame_vm_group_bin_11040 (RW)
0x68: frame_vm_group_bin_3855 (RW)
0x69: frame_vm_group_bin_19953 (RW)
0x6: frame_vm_group_bin_7131 (RW)
0x6a: frame_vm_group_bin_12752 (RW)
0x6b: frame_vm_group_bin_5688 (RW)
0x6c: frame_vm_group_bin_21787 (RW)
0x6d: frame_vm_group_bin_14613 (RW)
0x6e: frame_vm_group_bin_7399 (RW)
0x6f: frame_vm_group_bin_3940 (RW)
0x70: frame_vm_group_bin_16428 (RW)
0x71: frame_vm_group_bin_9238 (RW)
0x72: frame_vm_group_bin_2065 (RW)
0x73: frame_vm_group_bin_18161 (RW)
0x74: frame_vm_group_bin_11073 (RW)
0x75: frame_vm_group_bin_3888 (RW)
0x76: frame_vm_group_bin_19986 (RW)
0x77: frame_vm_group_bin_12785 (RW)
0x78: frame_vm_group_bin_5721 (RW)
0x79: frame_vm_group_bin_21821 (RW)
0x7: frame_vm_group_bin_0052 (RW)
0x7a: frame_vm_group_bin_14647 (RW)
0x7b: frame_vm_group_bin_7433 (RW)
0x7c: frame_vm_group_bin_8577 (RW)
0x7d: frame_vm_group_bin_16462 (RW)
0x7e: frame_vm_group_bin_9262 (RW)
0x7f: frame_vm_group_bin_2099 (RW)
0x80: frame_vm_group_bin_18194 (RW)
0x81: frame_vm_group_bin_11107 (RW)
0x82: frame_vm_group_bin_3922 (RW)
0x83: frame_vm_group_bin_20018 (RW)
0x84: frame_vm_group_bin_12818 (RW)
0x85: frame_vm_group_bin_5751 (RW)
0x86: frame_vm_group_bin_21855 (RW)
0x87: frame_vm_group_bin_14680 (RW)
0x88: frame_vm_group_bin_7466 (RW)
0x89: frame_vm_group_bin_0313 (RW)
0x8: frame_vm_group_bin_16180 (RW)
0x8a: frame_vm_group_bin_16495 (RW)
0x8b: frame_vm_group_bin_9287 (RW)
0x8c: frame_vm_group_bin_2133 (RW)
0x8d: frame_vm_group_bin_18227 (RW)
0x8e: frame_vm_group_bin_11139 (RW)
0x8f: frame_vm_group_bin_3954 (RW)
0x90: frame_vm_group_bin_20051 (RW)
0x91: frame_vm_group_bin_12851 (RW)
0x92: frame_vm_group_bin_5774 (RW)
0x93: frame_vm_group_bin_21888 (RW)
0x94: frame_vm_group_bin_14713 (RW)
0x95: frame_vm_group_bin_7499 (RW)
0x96: frame_vm_group_bin_17870 (RW)
0x97: frame_vm_group_bin_16528 (RW)
0x98: frame_vm_group_bin_9316 (RW)
0x99: frame_vm_group_bin_2166 (RW)
0x9: frame_vm_group_bin_8987 (RW)
0x9a: frame_vm_group_bin_18261 (RW)
0x9b: frame_vm_group_bin_11173 (RW)
0x9c: frame_vm_group_bin_3988 (RW)
0x9d: frame_vm_group_bin_20085 (RW)
0x9e: frame_vm_group_bin_12885 (RW)
0x9f: frame_vm_group_bin_22526 (RW)
0xa0: frame_vm_group_bin_21921 (RW)
0xa1: frame_vm_group_bin_14746 (RW)
0xa2: frame_vm_group_bin_7531 (RW)
0xa3: frame_vm_group_bin_0377 (RW)
0xa4: frame_vm_group_bin_16561 (RW)
0xa5: frame_vm_group_bin_9350 (RW)
0xa6: frame_vm_group_bin_2199 (RW)
0xa7: frame_vm_group_bin_18294 (RW)
0xa8: frame_vm_group_bin_11206 (RW)
0xa9: frame_vm_group_bin_4021 (RW)
0xa: frame_vm_group_bin_1799 (RW)
0xaa: frame_vm_group_bin_20117 (RW)
0xab: frame_vm_group_bin_12918 (RW)
0xac: frame_vm_group_bin_9675 (RW)
0xad: frame_vm_group_bin_21954 (RW)
0xae: frame_vm_group_bin_14778 (RW)
0xaf: frame_vm_group_bin_7563 (RW)
0xb0: frame_vm_group_bin_3962 (RW)
0xb1: frame_vm_group_bin_16594 (RW)
0xb2: frame_vm_group_bin_9383 (RW)
0xb3: frame_vm_group_bin_2228 (RW)
0xb4: frame_vm_group_bin_18327 (RW)
0xb5: frame_vm_group_bin_11239 (RW)
0xb6: frame_vm_group_bin_4054 (RW)
0xb7: frame_vm_group_bin_20150 (RW)
0xb8: frame_vm_group_bin_12950 (RW)
0xb9: frame_vm_group_bin_14338 (RW)
0xb: frame_vm_group_bin_17902 (RW)
0xba: frame_vm_group_bin_21988 (RW)
0xbb: frame_vm_group_bin_14812 (RW)
0xbc: frame_vm_group_bin_7597 (RW)
0xbd: frame_vm_group_bin_0437 (RW)
0xbe: frame_vm_group_bin_16627 (RW)
0xbf: frame_vm_group_bin_9418 (RW)
0xc0: frame_vm_group_bin_2258 (RW)
0xc1: frame_vm_group_bin_18361 (RW)
0xc2: frame_vm_group_bin_11273 (RW)
0xc3: frame_vm_group_bin_4088 (RW)
0xc4: frame_vm_group_bin_20182 (RW)
0xc5: frame_vm_group_bin_12984 (RW)
0xc6: frame_vm_group_bin_18964 (RW)
0xc7: frame_vm_group_bin_22019 (RW)
0xc8: frame_vm_group_bin_14845 (RW)
0xc9: frame_vm_group_bin_7630 (RW)
0xc: frame_vm_group_bin_10807 (RW)
0xca: frame_vm_group_bin_0470 (RW)
0xcb: frame_vm_group_bin_16660 (RW)
0xcc: frame_vm_group_bin_9451 (RW)
0xcd: frame_vm_group_bin_2291 (RW)
0xce: frame_vm_group_bin_18393 (RW)
0xcf: frame_vm_group_bin_11306 (RW)
0xd0: frame_vm_group_bin_4120 (RW)
0xd1: frame_vm_group_bin_20215 (RW)
0xd2: frame_vm_group_bin_13019 (RW)
0xd3: frame_vm_group_bin_5893 (RW)
0xd4: frame_vm_group_bin_22042 (RW)
0xd5: frame_vm_group_bin_14878 (RW)
0xd6: frame_vm_group_bin_7663 (RW)
0xd7: frame_vm_group_bin_0502 (RW)
0xd8: frame_vm_group_bin_16693 (RW)
0xd9: frame_vm_group_bin_9484 (RW)
0xd: frame_vm_group_bin_3622 (RW)
0xda: frame_vm_group_bin_2325 (RW)
0xdb: frame_vm_group_bin_18426 (RW)
0xdc: frame_vm_group_bin_11340 (RW)
0xdd: frame_vm_group_bin_4154 (RW)
0xde: frame_vm_group_bin_20249 (RW)
0xdf: frame_vm_group_bin_13053 (RW)
0xe0: frame_vm_group_bin_5070 (RW)
0xe1: frame_vm_group_bin_22067 (RW)
0xe2: frame_vm_group_bin_14912 (RW)
0xe3: frame_vm_group_bin_7697 (RW)
0xe4: frame_vm_group_bin_0535 (RW)
0xe5: frame_vm_group_bin_16727 (RW)
0xe6: frame_vm_group_bin_9518 (RW)
0xe7: frame_vm_group_bin_2358 (RW)
0xe8: frame_vm_group_bin_18458 (RW)
0xe9: frame_vm_group_bin_11371 (RW)
0xe: frame_vm_group_bin_19722 (RW)
0xea: frame_vm_group_bin_4186 (RW)
0xeb: frame_vm_group_bin_20281 (RW)
0xec: frame_vm_group_bin_13086 (RW)
0xed: frame_vm_group_bin_9699 (RW)
0xee: frame_vm_group_bin_22095 (RW)
0xef: frame_vm_group_bin_14945 (RW)
0xf0: frame_vm_group_bin_7729 (RW)
0xf1: frame_vm_group_bin_0566 (RW)
0xf2: frame_vm_group_bin_16760 (RW)
0xf3: frame_vm_group_bin_9551 (RW)
0xf4: frame_vm_group_bin_2391 (RW)
0xf5: frame_vm_group_bin_18485 (RW)
0xf6: frame_vm_group_bin_11403 (RW)
0xf7: frame_vm_group_bin_4218 (RW)
0xf8: frame_vm_group_bin_20314 (RW)
0xf9: frame_vm_group_bin_13119 (RW)
0xf: frame_vm_group_bin_12550 (RW)
0xfa: frame_vm_group_bin_14361 (RW)
0xfb: frame_vm_group_bin_22128 (RW)
0xfc: frame_vm_group_bin_14979 (RW)
0xfd: frame_vm_group_bin_7763 (RW)
0xfe: frame_vm_group_bin_0599 (RW)
0xff: frame_vm_group_bin_16794 (RW)
}
pt_vm_group_bin_0099 {
0x0: frame_vm_group_bin_13383 (RW)
0x100: frame_vm_group_bin_19393 (RW)
0x101: frame_vm_group_bin_12212 (RW)
0x102: frame_vm_group_bin_5122 (RW)
0x103: frame_vm_group_bin_21218 (RW)
0x104: frame_vm_group_bin_14041 (RW)
0x105: frame_vm_group_bin_6852 (RW)
0x106: frame_vm_group_bin_23055 (RW)
0x107: frame_vm_group_bin_15872 (RW)
0x108: frame_vm_group_bin_5935 (RW)
0x109: frame_vm_group_bin_1492 (RW)
0x10: frame_vm_group_bin_15242 (RW)
0x10a: frame_vm_group_bin_17632 (RW)
0x10b: frame_vm_group_bin_10503 (RW)
0x10c: frame_vm_group_bin_3356 (RW)
0x10d: frame_vm_group_bin_19425 (RW)
0x10e: frame_vm_group_bin_12244 (RW)
0x10f: frame_vm_group_bin_5155 (RW)
0x110: frame_vm_group_bin_21251 (RW)
0x111: frame_vm_group_bin_14074 (RW)
0x112: frame_vm_group_bin_6877 (RW)
0x113: frame_vm_group_bin_23088 (RW)
0x114: frame_vm_group_bin_15905 (RW)
0x115: frame_vm_group_bin_8714 (RW)
0x116: frame_vm_group_bin_1525 (RW)
0x117: frame_vm_group_bin_17665 (RW)
0x118: frame_vm_group_bin_10535 (RW)
0x119: frame_vm_group_bin_3386 (RW)
0x11: frame_vm_group_bin_8053 (RW)
0x11a: frame_vm_group_bin_19456 (RW)
0x11b: frame_vm_group_bin_2000 (RW)
0x11c: frame_vm_group_bin_5189 (RW)
0x11d: frame_vm_group_bin_21285 (RW)
0x11e: frame_vm_group_bin_14108 (RW)
0x11f: frame_vm_group_bin_6902 (RW)
0x120: frame_vm_group_bin_23122 (RW)
0x121: frame_vm_group_bin_15939 (RW)
0x122: frame_vm_group_bin_8748 (RW)
0x123: frame_vm_group_bin_1559 (RW)
0x124: frame_vm_group_bin_17695 (RW)
0x125: frame_vm_group_bin_10569 (RW)
0x126: frame_vm_group_bin_3414 (RW)
0x127: frame_vm_group_bin_19489 (RW)
0x128: frame_vm_group_bin_12311 (RW)
0x129: frame_vm_group_bin_5222 (RW)
0x12: frame_vm_group_bin_0896 (RW)
0x12a: frame_vm_group_bin_21317 (RW)
0x12b: frame_vm_group_bin_14141 (RW)
0x12c: frame_vm_group_bin_6930 (RW)
0x12d: frame_vm_group_bin_23154 (RW)
0x12e: frame_vm_group_bin_15972 (RW)
0x12f: frame_vm_group_bin_8781 (RW)
0x130: frame_vm_group_bin_1592 (RW)
0x131: frame_vm_group_bin_17122 (RW)
0x132: frame_vm_group_bin_10602 (RW)
0x133: frame_vm_group_bin_3436 (RW)
0x134: frame_vm_group_bin_19522 (RW)
0x135: frame_vm_group_bin_12343 (RW)
0x136: frame_vm_group_bin_5255 (RW)
0x137: frame_vm_group_bin_21349 (RW)
0x138: frame_vm_group_bin_14174 (RW)
0x139: frame_vm_group_bin_6961 (RW)
0x13: frame_vm_group_bin_17091 (RW)
0x13a: frame_vm_group_bin_23187 (RW)
0x13b: frame_vm_group_bin_16008 (RW)
0x13c: frame_vm_group_bin_8815 (RW)
0x13d: frame_vm_group_bin_1626 (RW)
0x13e: frame_vm_group_bin_17748 (RW)
0x13f: frame_vm_group_bin_10636 (RW)
0x140: frame_vm_group_bin_3462 (RW)
0x141: frame_vm_group_bin_19556 (RW)
0x142: frame_vm_group_bin_12377 (RW)
0x143: frame_vm_group_bin_5289 (RW)
0x144: frame_vm_group_bin_21383 (RW)
0x145: frame_vm_group_bin_14207 (RW)
0x146: frame_vm_group_bin_6994 (RW)
0x147: frame_vm_group_bin_23214 (RW)
0x148: frame_vm_group_bin_16041 (RW)
0x149: frame_vm_group_bin_8848 (RW)
0x14: frame_vm_group_bin_9883 (RW)
0x14a: frame_vm_group_bin_1659 (RW)
0x14b: frame_vm_group_bin_17778 (RW)
0x14c: frame_vm_group_bin_10667 (RW)
0x14d: frame_vm_group_bin_3488 (RW)
0x14e: frame_vm_group_bin_19590 (RW)
0x14f: frame_vm_group_bin_12410 (RW)
0x150: frame_vm_group_bin_5321 (RW)
0x151: frame_vm_group_bin_21416 (RW)
0x152: frame_vm_group_bin_14240 (RW)
0x153: frame_vm_group_bin_7027 (RW)
0x154: frame_vm_group_bin_23236 (RW)
0x155: frame_vm_group_bin_16074 (RW)
0x156: frame_vm_group_bin_8880 (RW)
0x157: frame_vm_group_bin_1692 (RW)
0x158: frame_vm_group_bin_17809 (RW)
0x159: frame_vm_group_bin_10700 (RW)
0x15: frame_vm_group_bin_2722 (RW)
0x15a: frame_vm_group_bin_3516 (RW)
0x15b: frame_vm_group_bin_19624 (RW)
0x15c: frame_vm_group_bin_12443 (RW)
0x15d: frame_vm_group_bin_5353 (RW)
0x15e: frame_vm_group_bin_21449 (RW)
0x15f: frame_vm_group_bin_14273 (RW)
0x160: frame_vm_group_bin_7059 (RW)
0x161: frame_vm_group_bin_0641 (RW)
0x162: frame_vm_group_bin_16107 (RW)
0x163: frame_vm_group_bin_8913 (RW)
0x164: frame_vm_group_bin_1725 (RW)
0x165: frame_vm_group_bin_17838 (RW)
0x166: frame_vm_group_bin_10733 (RW)
0x167: frame_vm_group_bin_3547 (RW)
0x168: frame_vm_group_bin_19654 (RW)
0x169: frame_vm_group_bin_12475 (RW)
0x16: frame_vm_group_bin_18795 (RW)
0x16a: frame_vm_group_bin_5385 (RW)
0x16b: frame_vm_group_bin_21481 (RW)
0x16c: frame_vm_group_bin_14304 (RW)
0x16d: frame_vm_group_bin_7091 (RW)
0x16e: frame_vm_group_bin_22858 (RW)
0x16f: frame_vm_group_bin_16138 (RW)
0x170: frame_vm_group_bin_8945 (RW)
0x171: frame_vm_group_bin_1757 (RW)
0x172: frame_vm_group_bin_17145 (RW)
0x173: frame_vm_group_bin_10766 (RW)
0x174: frame_vm_group_bin_3579 (RW)
0x175: frame_vm_group_bin_19681 (RW)
0x176: frame_vm_group_bin_12508 (RW)
0x177: frame_vm_group_bin_5418 (RW)
0x178: frame_vm_group_bin_21513 (RW)
0x179: frame_vm_group_bin_14337 (RW)
0x17: frame_vm_group_bin_1906 (RW)
0x17a: frame_vm_group_bin_7124 (RW)
0x17b: frame_vm_group_bin_4221 (RW)
0x17c: frame_vm_group_bin_16172 (RW)
0x17d: frame_vm_group_bin_8979 (RW)
0x17e: frame_vm_group_bin_1791 (RW)
0x17f: frame_vm_group_bin_21776 (RW)
0x180: frame_vm_group_bin_10799 (RW)
0x181: frame_vm_group_bin_3614 (RW)
0x182: frame_vm_group_bin_19714 (RW)
0x183: frame_vm_group_bin_12542 (RW)
0x184: frame_vm_group_bin_5451 (RW)
0x185: frame_vm_group_bin_21547 (RW)
0x186: frame_vm_group_bin_14371 (RW)
0x187: frame_vm_group_bin_7156 (RW)
0x188: frame_vm_group_bin_0071 (RW)
0x189: frame_vm_group_bin_16203 (RW)
0x18: frame_vm_group_bin_4552 (RW)
0x18a: frame_vm_group_bin_9012 (RW)
0x18b: frame_vm_group_bin_1824 (RW)
0x18c: frame_vm_group_bin_17926 (RW)
0x18d: frame_vm_group_bin_10832 (RW)
0x18e: frame_vm_group_bin_3647 (RW)
0x18f: frame_vm_group_bin_19747 (RW)
0x190: frame_vm_group_bin_12575 (RW)
0x191: frame_vm_group_bin_5483 (RW)
0x192: frame_vm_group_bin_21580 (RW)
0x193: frame_vm_group_bin_14404 (RW)
0x194: frame_vm_group_bin_7191 (RW)
0x195: frame_vm_group_bin_13499 (RW)
0x196: frame_vm_group_bin_16230 (RW)
0x197: frame_vm_group_bin_9045 (RW)
0x198: frame_vm_group_bin_1857 (RW)
0x199: frame_vm_group_bin_17957 (RW)
0x19: frame_vm_group_bin_20649 (RW)
0x19a: frame_vm_group_bin_10866 (RW)
0x19b: frame_vm_group_bin_3681 (RW)
0x19c: frame_vm_group_bin_19781 (RW)
0x19d: frame_vm_group_bin_12609 (RW)
0x19e: frame_vm_group_bin_5516 (RW)
0x19f: frame_vm_group_bin_21614 (RW)
0x1: frame_vm_group_bin_10174 (RW)
0x1a0: frame_vm_group_bin_14438 (RW)
0x1a1: frame_vm_group_bin_7225 (RW)
0x1a2: frame_vm_group_bin_18143 (RW)
0x1a3: frame_vm_group_bin_16259 (RW)
0x1a4: frame_vm_group_bin_9079 (RW)
0x1a5: frame_vm_group_bin_1891 (RW)
0x1a6: frame_vm_group_bin_17989 (RW)
0x1a7: frame_vm_group_bin_10899 (RW)
0x1a8: frame_vm_group_bin_3714 (RW)
0x1a9: frame_vm_group_bin_19814 (RW)
0x1a: frame_vm_group_bin_13450 (RW)
0x1aa: frame_vm_group_bin_12641 (RW)
0x1ab: frame_vm_group_bin_5549 (RW)
0x1ac: frame_vm_group_bin_21647 (RW)
0x1ad: frame_vm_group_bin_14471 (RW)
0x1ae: frame_vm_group_bin_7258 (RW)
0x1af: frame_vm_group_bin_22882 (RW)
0x1b0: frame_vm_group_bin_16288 (RW)
0x1b1: frame_vm_group_bin_9112 (RW)
0x1b2: frame_vm_group_bin_1924 (RW)
0x1b3: frame_vm_group_bin_18022 (RW)
0x1b4: frame_vm_group_bin_10932 (RW)
0x1b5: frame_vm_group_bin_3747 (RW)
0x1b6: frame_vm_group_bin_19847 (RW)
0x1b7: frame_vm_group_bin_12668 (RW)
0x1b8: frame_vm_group_bin_5581 (RW)
0x1b9: frame_vm_group_bin_21679 (RW)
0x1b: frame_vm_group_bin_19455 (RW)
0x1ba: frame_vm_group_bin_14506 (RW)
0x1bb: frame_vm_group_bin_7291 (RW)
0x1bc: frame_vm_group_bin_0167 (RW)
0x1bd: frame_vm_group_bin_16320 (RW)
0x1be: frame_vm_group_bin_9145 (RW)
0x1bf: frame_vm_group_bin_1957 (RW)
0x1c0: frame_vm_group_bin_18055 (RW)
0x1c1: frame_vm_group_bin_10965 (RW)
0x1c2: frame_vm_group_bin_3780 (RW)
0x1c3: frame_vm_group_bin_19880 (RW)
0x1c4: frame_vm_group_bin_12694 (RW)
0x1c5: frame_vm_group_bin_5613 (RW)
0x1c6: frame_vm_group_bin_21713 (RW)
0x1c7: frame_vm_group_bin_14539 (RW)
0x1c8: frame_vm_group_bin_7324 (RW)
0x1c9: frame_vm_group_bin_0198 (RW)
0x1c: frame_vm_group_bin_22458 (RW)
0x1ca: frame_vm_group_bin_16353 (RW)
0x1cb: frame_vm_group_bin_9177 (RW)
0x1cc: frame_vm_group_bin_1990 (RW)
0x1cd: frame_vm_group_bin_18087 (RW)
0x1ce: frame_vm_group_bin_10998 (RW)
0x1cf: frame_vm_group_bin_3813 (RW)
0x1d0: frame_vm_group_bin_19912 (RW)
0x1d1: frame_vm_group_bin_12719 (RW)
0x1d2: frame_vm_group_bin_5646 (RW)
0x1d3: frame_vm_group_bin_21746 (RW)
0x1d4: frame_vm_group_bin_14572 (RW)
0x1d5: frame_vm_group_bin_7357 (RW)
0x1d6: frame_vm_group_bin_0228 (RW)
0x1d7: frame_vm_group_bin_16386 (RW)
0x1d8: frame_vm_group_bin_9205 (RW)
0x1d9: frame_vm_group_bin_2023 (RW)
0x1d: frame_vm_group_bin_15276 (RW)
0x1da: frame_vm_group_bin_18120 (RW)
0x1db: frame_vm_group_bin_11032 (RW)
0x1dc: frame_vm_group_bin_3847 (RW)
0x1dd: frame_vm_group_bin_19945 (RW)
0x1de: frame_vm_group_bin_12745 (RW)
0x1df: frame_vm_group_bin_5680 (RW)
0x1e0: frame_vm_group_bin_21779 (RW)
0x1e1: frame_vm_group_bin_14605 (RW)
0x1e2: frame_vm_group_bin_7391 (RW)
0x1e3: frame_vm_group_bin_18168 (RW)
0x1e4: frame_vm_group_bin_16420 (RW)
0x1e5: frame_vm_group_bin_9233 (RW)
0x1e6: frame_vm_group_bin_2057 (RW)
0x1e7: frame_vm_group_bin_18153 (RW)
0x1e8: frame_vm_group_bin_11065 (RW)
0x1e9: frame_vm_group_bin_3880 (RW)
0x1e: frame_vm_group_bin_8085 (RW)
0x1ea: frame_vm_group_bin_19978 (RW)
0x1eb: frame_vm_group_bin_12777 (RW)
0x1ec: frame_vm_group_bin_5713 (RW)
0x1ed: frame_vm_group_bin_21813 (RW)
0x1ee: frame_vm_group_bin_14638 (RW)
0x1ef: frame_vm_group_bin_7424 (RW)
0x1f0: frame_vm_group_bin_0275 (RW)
0x1f1: frame_vm_group_bin_16453 (RW)
0x1f2: frame_vm_group_bin_9256 (RW)
0x1f3: frame_vm_group_bin_2090 (RW)
0x1f4: frame_vm_group_bin_18186 (RW)
0x1f5: frame_vm_group_bin_11098 (RW)
0x1f6: frame_vm_group_bin_3913 (RW)
0x1f7: frame_vm_group_bin_20009 (RW)
0x1f8: frame_vm_group_bin_12810 (RW)
0x1f9: frame_vm_group_bin_5743 (RW)
0x1f: frame_vm_group_bin_0930 (RW)
0x1fa: frame_vm_group_bin_21847 (RW)
0x1fb: frame_vm_group_bin_14672 (RW)
0x1fc: frame_vm_group_bin_7458 (RW)
0x1fd: frame_vm_group_bin_0305 (RW)
0x1fe: frame_vm_group_bin_16487 (RW)
0x1ff: frame_vm_group_bin_9282 (RW)
0x20: frame_vm_group_bin_17125 (RW)
0x21: frame_vm_group_bin_9916 (RW)
0x22: frame_vm_group_bin_2756 (RW)
0x23: frame_vm_group_bin_18830 (RW)
0x24: frame_vm_group_bin_6544 (RW)
0x25: frame_vm_group_bin_4581 (RW)
0x26: frame_vm_group_bin_20682 (RW)
0x27: frame_vm_group_bin_13483 (RW)
0x28: frame_vm_group_bin_6298 (RW)
0x29: frame_vm_group_bin_22491 (RW)
0x2: frame_vm_group_bin_22392 (RW)
0x2a: frame_vm_group_bin_15308 (RW)
0x2b: frame_vm_group_bin_8117 (RW)
0x2c: frame_vm_group_bin_0963 (RW)
0x2d: frame_vm_group_bin_17157 (RW)
0x2e: frame_vm_group_bin_9947 (RW)
0x2f: frame_vm_group_bin_2789 (RW)
0x30: frame_vm_group_bin_18863 (RW)
0x31: frame_vm_group_bin_11291 (RW)
0x32: frame_vm_group_bin_4603 (RW)
0x33: frame_vm_group_bin_20715 (RW)
0x34: frame_vm_group_bin_13516 (RW)
0x35: frame_vm_group_bin_6330 (RW)
0x36: frame_vm_group_bin_22524 (RW)
0x37: frame_vm_group_bin_15341 (RW)
0x38: frame_vm_group_bin_8150 (RW)
0x39: frame_vm_group_bin_0996 (RW)
0x3: frame_vm_group_bin_15208 (RW)
0x3a: frame_vm_group_bin_17190 (RW)
0x3b: frame_vm_group_bin_9981 (RW)
0x3c: frame_vm_group_bin_2823 (RW)
0x3d: frame_vm_group_bin_18897 (RW)
0x3e: frame_vm_group_bin_11763 (RW)
0x3f: frame_vm_group_bin_4629 (RW)
0x40: frame_vm_group_bin_20749 (RW)
0x41: frame_vm_group_bin_13550 (RW)
0x42: frame_vm_group_bin_6364 (RW)
0x43: frame_vm_group_bin_22557 (RW)
0x44: frame_vm_group_bin_15375 (RW)
0x45: frame_vm_group_bin_8184 (RW)
0x46: frame_vm_group_bin_1025 (RW)
0x47: frame_vm_group_bin_17221 (RW)
0x48: frame_vm_group_bin_10014 (RW)
0x49: frame_vm_group_bin_0149 (RW)
0x4: frame_vm_group_bin_5862 (RW)
0x4a: frame_vm_group_bin_18930 (RW)
0x4b: frame_vm_group_bin_20581 (RW)
0x4c: frame_vm_group_bin_4661 (RW)
0x4d: frame_vm_group_bin_20782 (RW)
0x4e: frame_vm_group_bin_13583 (RW)
0x4f: frame_vm_group_bin_6394 (RW)
0x50: frame_vm_group_bin_22590 (RW)
0x51: frame_vm_group_bin_15408 (RW)
0x52: frame_vm_group_bin_8217 (RW)
0x53: frame_vm_group_bin_1047 (RW)
0x54: frame_vm_group_bin_17253 (RW)
0x55: frame_vm_group_bin_10047 (RW)
0x56: frame_vm_group_bin_2890 (RW)
0x57: frame_vm_group_bin_18962 (RW)
0x58: frame_vm_group_bin_11819 (RW)
0x59: frame_vm_group_bin_4693 (RW)
0x5: frame_vm_group_bin_0863 (RW)
0x5a: frame_vm_group_bin_20816 (RW)
0x5b: frame_vm_group_bin_13617 (RW)
0x5c: frame_vm_group_bin_6427 (RW)
0x5d: frame_vm_group_bin_22624 (RW)
0x5e: frame_vm_group_bin_15442 (RW)
0x5f: frame_vm_group_bin_8251 (RW)
0x60: frame_vm_group_bin_1071 (RW)
0x61: frame_vm_group_bin_17287 (RW)
0x62: frame_vm_group_bin_10081 (RW)
0x63: frame_vm_group_bin_2924 (RW)
0x64: frame_vm_group_bin_18994 (RW)
0x65: frame_vm_group_bin_11850 (RW)
0x66: frame_vm_group_bin_4725 (RW)
0x67: frame_vm_group_bin_20846 (RW)
0x68: frame_vm_group_bin_13649 (RW)
0x69: frame_vm_group_bin_6460 (RW)
0x6: frame_vm_group_bin_17058 (RW)
0x6a: frame_vm_group_bin_22657 (RW)
0x6b: frame_vm_group_bin_15475 (RW)
0x6c: frame_vm_group_bin_8283 (RW)
0x6d: frame_vm_group_bin_1097 (RW)
0x6e: frame_vm_group_bin_17320 (RW)
0x6f: frame_vm_group_bin_10114 (RW)
0x70: frame_vm_group_bin_2957 (RW)
0x71: frame_vm_group_bin_19027 (RW)
0x72: frame_vm_group_bin_11879 (RW)
0x73: frame_vm_group_bin_4758 (RW)
0x74: frame_vm_group_bin_20870 (RW)
0x75: frame_vm_group_bin_13682 (RW)
0x76: frame_vm_group_bin_6493 (RW)
0x77: frame_vm_group_bin_22690 (RW)
0x78: frame_vm_group_bin_15508 (RW)
0x79: frame_vm_group_bin_8316 (RW)
0x7: frame_vm_group_bin_9850 (RW)
0x7a: frame_vm_group_bin_1128 (RW)
0x7b: frame_vm_group_bin_17354 (RW)
0x7c: frame_vm_group_bin_10150 (RW)
0x7d: frame_vm_group_bin_2991 (RW)
0x7e: frame_vm_group_bin_19061 (RW)
0x7f: frame_vm_group_bin_11903 (RW)
0x80: frame_vm_group_bin_4792 (RW)
0x81: frame_vm_group_bin_20900 (RW)
0x82: frame_vm_group_bin_13715 (RW)
0x83: frame_vm_group_bin_6527 (RW)
0x84: frame_vm_group_bin_22724 (RW)
0x85: frame_vm_group_bin_15540 (RW)
0x86: frame_vm_group_bin_8350 (RW)
0x87: frame_vm_group_bin_1161 (RW)
0x88: frame_vm_group_bin_17385 (RW)
0x89: frame_vm_group_bin_10183 (RW)
0x8: frame_vm_group_bin_2689 (RW)
0x8a: frame_vm_group_bin_3024 (RW)
0x8b: frame_vm_group_bin_19094 (RW)
0x8c: frame_vm_group_bin_11932 (RW)
0x8d: frame_vm_group_bin_4824 (RW)
0x8e: frame_vm_group_bin_20925 (RW)
0x8f: frame_vm_group_bin_13748 (RW)
0x90: frame_vm_group_bin_6560 (RW)
0x91: frame_vm_group_bin_22756 (RW)
0x92: frame_vm_group_bin_15573 (RW)
0x93: frame_vm_group_bin_8383 (RW)
0x94: frame_vm_group_bin_1194 (RW)
0x95: frame_vm_group_bin_17411 (RW)
0x96: frame_vm_group_bin_10216 (RW)
0x97: frame_vm_group_bin_3057 (RW)
0x98: frame_vm_group_bin_19126 (RW)
0x99: frame_vm_group_bin_11962 (RW)
0x9: frame_vm_group_bin_18762 (RW)
0x9a: frame_vm_group_bin_4858 (RW)
0x9b: frame_vm_group_bin_20953 (RW)
0x9c: frame_vm_group_bin_13783 (RW)
0x9d: frame_vm_group_bin_6594 (RW)
0x9e: frame_vm_group_bin_22790 (RW)
0x9f: frame_vm_group_bin_15607 (RW)
0xa0: frame_vm_group_bin_8417 (RW)
0xa1: frame_vm_group_bin_1228 (RW)
0xa2: frame_vm_group_bin_17439 (RW)
0xa3: frame_vm_group_bin_10250 (RW)
0xa4: frame_vm_group_bin_3091 (RW)
0xa5: frame_vm_group_bin_19159 (RW)
0xa6: frame_vm_group_bin_11995 (RW)
0xa7: frame_vm_group_bin_4891 (RW)
0xa8: frame_vm_group_bin_20984 (RW)
0xa9: frame_vm_group_bin_13815 (RW)
0xa: frame_vm_group_bin_20557 (RW)
0xaa: frame_vm_group_bin_6627 (RW)
0xab: frame_vm_group_bin_22823 (RW)
0xac: frame_vm_group_bin_15640 (RW)
0xad: frame_vm_group_bin_8450 (RW)
0xae: frame_vm_group_bin_1260 (RW)
0xaf: frame_vm_group_bin_10888 (RW)
0xb0: frame_vm_group_bin_10283 (RW)
0xb1: frame_vm_group_bin_3123 (RW)
0xb2: frame_vm_group_bin_19192 (RW)
0xb3: frame_vm_group_bin_12026 (RW)
0xb4: frame_vm_group_bin_4923 (RW)
0xb5: frame_vm_group_bin_21017 (RW)
0xb6: frame_vm_group_bin_13844 (RW)
0xb7: frame_vm_group_bin_6660 (RW)
0xb8: frame_vm_group_bin_22856 (RW)
0xb9: frame_vm_group_bin_15673 (RW)
0xb: frame_vm_group_bin_4520 (RW)
0xba: frame_vm_group_bin_8484 (RW)
0xbb: frame_vm_group_bin_1292 (RW)
0xbc: frame_vm_group_bin_21703 (RW)
0xbd: frame_vm_group_bin_10317 (RW)
0xbe: frame_vm_group_bin_3157 (RW)
0xbf: frame_vm_group_bin_19226 (RW)
0xc0: frame_vm_group_bin_15983 (RW)
0xc1: frame_vm_group_bin_4955 (RW)
0xc2: frame_vm_group_bin_21052 (RW)
0xc3: frame_vm_group_bin_13875 (RW)
0xc4: frame_vm_group_bin_6694 (RW)
0xc5: frame_vm_group_bin_22890 (RW)
0xc6: frame_vm_group_bin_15707 (RW)
0xc7: frame_vm_group_bin_8516 (RW)
0xc8: frame_vm_group_bin_1324 (RW)
0xc9: frame_vm_group_bin_3084 (RW)
0xc: frame_vm_group_bin_20616 (RW)
0xca: frame_vm_group_bin_10350 (RW)
0xcb: frame_vm_group_bin_3190 (RW)
0xcc: frame_vm_group_bin_19259 (RW)
0xcd: frame_vm_group_bin_12086 (RW)
0xce: frame_vm_group_bin_4987 (RW)
0xcf: frame_vm_group_bin_21085 (RW)
0xd0: frame_vm_group_bin_13907 (RW)
0xd1: frame_vm_group_bin_6726 (RW)
0xd2: frame_vm_group_bin_22923 (RW)
0xd3: frame_vm_group_bin_15740 (RW)
0xd4: frame_vm_group_bin_8548 (RW)
0xd5: frame_vm_group_bin_1357 (RW)
0xd6: frame_vm_group_bin_7691 (RW)
0xd7: frame_vm_group_bin_10382 (RW)
0xd8: frame_vm_group_bin_3223 (RW)
0xd9: frame_vm_group_bin_19292 (RW)
0xd: frame_vm_group_bin_13416 (RW)
0xda: frame_vm_group_bin_12119 (RW)
0xdb: frame_vm_group_bin_5021 (RW)
0xdc: frame_vm_group_bin_21119 (RW)
0xdd: frame_vm_group_bin_13941 (RW)
0xde: frame_vm_group_bin_6759 (RW)
0xdf: frame_vm_group_bin_22956 (RW)
0xe0: frame_vm_group_bin_15774 (RW)
0xe1: frame_vm_group_bin_8581 (RW)
0xe2: frame_vm_group_bin_1392 (RW)
0xe3: frame_vm_group_bin_12348 (RW)
0xe4: frame_vm_group_bin_10410 (RW)
0xe5: frame_vm_group_bin_3256 (RW)
0xe6: frame_vm_group_bin_19326 (RW)
0xe7: frame_vm_group_bin_12152 (RW)
0xe8: frame_vm_group_bin_5054 (RW)
0xe9: frame_vm_group_bin_21151 (RW)
0xe: frame_vm_group_bin_14835 (RW)
0xea: frame_vm_group_bin_13974 (RW)
0xeb: frame_vm_group_bin_6792 (RW)
0xec: frame_vm_group_bin_22989 (RW)
0xed: frame_vm_group_bin_15806 (RW)
0xee: frame_vm_group_bin_8613 (RW)
0xef: frame_vm_group_bin_1425 (RW)
0xf0: frame_vm_group_bin_17098 (RW)
0xf1: frame_vm_group_bin_10438 (RW)
0xf2: frame_vm_group_bin_3289 (RW)
0xf3: frame_vm_group_bin_19359 (RW)
0xf4: frame_vm_group_bin_12182 (RW)
0xf5: frame_vm_group_bin_5088 (RW)
0xf6: frame_vm_group_bin_21184 (RW)
0xf7: frame_vm_group_bin_14007 (RW)
0xf8: frame_vm_group_bin_6822 (RW)
0xf9: frame_vm_group_bin_23021 (RW)
0xf: frame_vm_group_bin_22424 (RW)
0xfa: frame_vm_group_bin_15839 (RW)
0xfb: frame_vm_group_bin_8647 (RW)
0xfc: frame_vm_group_bin_1459 (RW)
0xfd: frame_vm_group_bin_21728 (RW)
0xfe: frame_vm_group_bin_10470 (RW)
0xff: frame_vm_group_bin_3323 (RW)
}
pt_vm_group_bin_0107 {
0x0: frame_vm_group_bin_17102 (RW)
0x100: frame_vm_group_bin_23099 (RW)
0x101: frame_vm_group_bin_15916 (RW)
0x102: frame_vm_group_bin_8725 (RW)
0x103: frame_vm_group_bin_1536 (RW)
0x104: frame_vm_group_bin_17676 (RW)
0x105: frame_vm_group_bin_10546 (RW)
0x106: frame_vm_group_bin_3397 (RW)
0x107: frame_vm_group_bin_19466 (RW)
0x108: frame_vm_group_bin_12288 (RW)
0x109: frame_vm_group_bin_5199 (RW)
0x10: frame_vm_group_bin_18840 (RW)
0x10a: frame_vm_group_bin_21295 (RW)
0x10b: frame_vm_group_bin_14118 (RW)
0x10c: frame_vm_group_bin_6909 (RW)
0x10d: frame_vm_group_bin_23132 (RW)
0x10e: frame_vm_group_bin_15949 (RW)
0x10f: frame_vm_group_bin_8758 (RW)
0x110: frame_vm_group_bin_1569 (RW)
0x111: frame_vm_group_bin_16365 (RW)
0x112: frame_vm_group_bin_10579 (RW)
0x113: frame_vm_group_bin_3421 (RW)
0x114: frame_vm_group_bin_19499 (RW)
0x115: frame_vm_group_bin_12321 (RW)
0x116: frame_vm_group_bin_5232 (RW)
0x117: frame_vm_group_bin_21327 (RW)
0x118: frame_vm_group_bin_14151 (RW)
0x119: frame_vm_group_bin_6939 (RW)
0x11: frame_vm_group_bin_10537 (RW)
0x11a: frame_vm_group_bin_23165 (RW)
0x11b: frame_vm_group_bin_15985 (RW)
0x11c: frame_vm_group_bin_8792 (RW)
0x11d: frame_vm_group_bin_1603 (RW)
0x11e: frame_vm_group_bin_17730 (RW)
0x11f: frame_vm_group_bin_10613 (RW)
0x120: frame_vm_group_bin_3444 (RW)
0x121: frame_vm_group_bin_19533 (RW)
0x122: frame_vm_group_bin_12354 (RW)
0x123: frame_vm_group_bin_5266 (RW)
0x124: frame_vm_group_bin_21360 (RW)
0x125: frame_vm_group_bin_14184 (RW)
0x126: frame_vm_group_bin_6971 (RW)
0x127: frame_vm_group_bin_23197 (RW)
0x128: frame_vm_group_bin_16018 (RW)
0x129: frame_vm_group_bin_8825 (RW)
0x12: frame_vm_group_bin_4588 (RW)
0x12a: frame_vm_group_bin_1636 (RW)
0x12b: frame_vm_group_bin_17757 (RW)
0x12c: frame_vm_group_bin_10645 (RW)
0x12d: frame_vm_group_bin_3469 (RW)
0x12e: frame_vm_group_bin_19566 (RW)
0x12f: frame_vm_group_bin_12387 (RW)
0x130: frame_vm_group_bin_5299 (RW)
0x131: frame_vm_group_bin_21393 (RW)
0x132: frame_vm_group_bin_14217 (RW)
0x133: frame_vm_group_bin_7004 (RW)
0x134: frame_vm_group_bin_23221 (RW)
0x135: frame_vm_group_bin_16051 (RW)
0x136: frame_vm_group_bin_8858 (RW)
0x137: frame_vm_group_bin_1669 (RW)
0x138: frame_vm_group_bin_17787 (RW)
0x139: frame_vm_group_bin_10677 (RW)
0x13: frame_vm_group_bin_20692 (RW)
0x13a: frame_vm_group_bin_3496 (RW)
0x13b: frame_vm_group_bin_19601 (RW)
0x13c: frame_vm_group_bin_12421 (RW)
0x13d: frame_vm_group_bin_5331 (RW)
0x13e: frame_vm_group_bin_21426 (RW)
0x13f: frame_vm_group_bin_14250 (RW)
0x140: frame_vm_group_bin_7037 (RW)
0x141: frame_vm_group_bin_23243 (RW)
0x142: frame_vm_group_bin_16084 (RW)
0x143: frame_vm_group_bin_8890 (RW)
0x144: frame_vm_group_bin_1702 (RW)
0x145: frame_vm_group_bin_17817 (RW)
0x146: frame_vm_group_bin_10710 (RW)
0x147: frame_vm_group_bin_3524 (RW)
0x148: frame_vm_group_bin_19633 (RW)
0x149: frame_vm_group_bin_12452 (RW)
0x14: frame_vm_group_bin_13493 (RW)
0x14a: frame_vm_group_bin_5362 (RW)
0x14b: frame_vm_group_bin_21458 (RW)
0x14c: frame_vm_group_bin_14282 (RW)
0x14d: frame_vm_group_bin_7068 (RW)
0x14e: frame_vm_group_bin_22103 (RW)
0x14f: frame_vm_group_bin_16116 (RW)
0x150: frame_vm_group_bin_8922 (RW)
0x151: frame_vm_group_bin_1734 (RW)
0x152: frame_vm_group_bin_17845 (RW)
0x153: frame_vm_group_bin_10742 (RW)
0x154: frame_vm_group_bin_3556 (RW)
0x155: frame_vm_group_bin_19661 (RW)
0x156: frame_vm_group_bin_12484 (RW)
0x157: frame_vm_group_bin_5394 (RW)
0x158: frame_vm_group_bin_21490 (RW)
0x159: frame_vm_group_bin_14313 (RW)
0x15: frame_vm_group_bin_6308 (RW)
0x15a: frame_vm_group_bin_7101 (RW)
0x15b: frame_vm_group_bin_3478 (RW)
0x15c: frame_vm_group_bin_16148 (RW)
0x15d: frame_vm_group_bin_8955 (RW)
0x15e: frame_vm_group_bin_1767 (RW)
0x15f: frame_vm_group_bin_17872 (RW)
0x160: frame_vm_group_bin_10775 (RW)
0x161: frame_vm_group_bin_3590 (RW)
0x162: frame_vm_group_bin_19690 (RW)
0x163: frame_vm_group_bin_12518 (RW)
0x164: frame_vm_group_bin_5428 (RW)
0x165: frame_vm_group_bin_21523 (RW)
0x166: frame_vm_group_bin_14347 (RW)
0x167: frame_vm_group_bin_7132 (RW)
0x168: frame_vm_group_bin_8107 (RW)
0x169: frame_vm_group_bin_16181 (RW)
0x16: frame_vm_group_bin_22501 (RW)
0x16a: frame_vm_group_bin_8988 (RW)
0x16b: frame_vm_group_bin_1800 (RW)
0x16c: frame_vm_group_bin_17903 (RW)
0x16d: frame_vm_group_bin_10808 (RW)
0x16e: frame_vm_group_bin_3623 (RW)
0x16f: frame_vm_group_bin_19723 (RW)
0x170: frame_vm_group_bin_12551 (RW)
0x171: frame_vm_group_bin_5460 (RW)
0x172: frame_vm_group_bin_21556 (RW)
0x173: frame_vm_group_bin_14380 (RW)
0x174: frame_vm_group_bin_7165 (RW)
0x175: frame_vm_group_bin_0078 (RW)
0x176: frame_vm_group_bin_16211 (RW)
0x177: frame_vm_group_bin_9021 (RW)
0x178: frame_vm_group_bin_1833 (RW)
0x179: frame_vm_group_bin_7010 (RW)
0x17: frame_vm_group_bin_15318 (RW)
0x17a: frame_vm_group_bin_10842 (RW)
0x17b: frame_vm_group_bin_3657 (RW)
0x17c: frame_vm_group_bin_19757 (RW)
0x17d: frame_vm_group_bin_12585 (RW)
0x17e: frame_vm_group_bin_5493 (RW)
0x17f: frame_vm_group_bin_21590 (RW)
0x180: frame_vm_group_bin_14414 (RW)
0x181: frame_vm_group_bin_7201 (RW)
0x182: frame_vm_group_bin_0104 (RW)
0x183: frame_vm_group_bin_16240 (RW)
0x184: frame_vm_group_bin_9055 (RW)
0x185: frame_vm_group_bin_1867 (RW)
0x186: frame_vm_group_bin_17967 (RW)
0x187: frame_vm_group_bin_10874 (RW)
0x188: frame_vm_group_bin_3690 (RW)
0x189: frame_vm_group_bin_19790 (RW)
0x18: frame_vm_group_bin_8127 (RW)
0x18a: frame_vm_group_bin_12618 (RW)
0x18b: frame_vm_group_bin_5525 (RW)
0x18c: frame_vm_group_bin_21623 (RW)
0x18d: frame_vm_group_bin_14447 (RW)
0x18e: frame_vm_group_bin_7234 (RW)
0x18f: frame_vm_group_bin_22126 (RW)
0x190: frame_vm_group_bin_16266 (RW)
0x191: frame_vm_group_bin_9088 (RW)
0x192: frame_vm_group_bin_1900 (RW)
0x193: frame_vm_group_bin_17998 (RW)
0x194: frame_vm_group_bin_10908 (RW)
0x195: frame_vm_group_bin_3723 (RW)
0x196: frame_vm_group_bin_19823 (RW)
0x197: frame_vm_group_bin_12649 (RW)
0x198: frame_vm_group_bin_5558 (RW)
0x199: frame_vm_group_bin_21656 (RW)
0x19: frame_vm_group_bin_0973 (RW)
0x19a: frame_vm_group_bin_14481 (RW)
0x19b: frame_vm_group_bin_7268 (RW)
0x19c: frame_vm_group_bin_3495 (RW)
0x19d: frame_vm_group_bin_16297 (RW)
0x19e: frame_vm_group_bin_9122 (RW)
0x19f: frame_vm_group_bin_1934 (RW)
0x1: frame_vm_group_bin_9893 (RW)
0x1a0: frame_vm_group_bin_18032 (RW)
0x1a1: frame_vm_group_bin_10942 (RW)
0x1a2: frame_vm_group_bin_3757 (RW)
0x1a3: frame_vm_group_bin_19857 (RW)
0x1a4: frame_vm_group_bin_12677 (RW)
0x1a5: frame_vm_group_bin_5591 (RW)
0x1a6: frame_vm_group_bin_21689 (RW)
0x1a7: frame_vm_group_bin_14515 (RW)
0x1a8: frame_vm_group_bin_7300 (RW)
0x1a9: frame_vm_group_bin_0175 (RW)
0x1a: frame_vm_group_bin_17168 (RW)
0x1aa: frame_vm_group_bin_16329 (RW)
0x1ab: frame_vm_group_bin_9154 (RW)
0x1ac: frame_vm_group_bin_1966 (RW)
0x1ad: frame_vm_group_bin_18064 (RW)
0x1ae: frame_vm_group_bin_10974 (RW)
0x1af: frame_vm_group_bin_3789 (RW)
0x1b0: frame_vm_group_bin_19889 (RW)
0x1b1: frame_vm_group_bin_12700 (RW)
0x1b2: frame_vm_group_bin_5622 (RW)
0x1b3: frame_vm_group_bin_21722 (RW)
0x1b4: frame_vm_group_bin_14548 (RW)
0x1b5: frame_vm_group_bin_7333 (RW)
0x1b6: frame_vm_group_bin_0207 (RW)
0x1b7: frame_vm_group_bin_16362 (RW)
0x1b8: frame_vm_group_bin_9185 (RW)
0x1b9: frame_vm_group_bin_1999 (RW)
0x1b: frame_vm_group_bin_9958 (RW)
0x1ba: frame_vm_group_bin_18098 (RW)
0x1bb: frame_vm_group_bin_11008 (RW)
0x1bc: frame_vm_group_bin_3823 (RW)
0x1bd: frame_vm_group_bin_19922 (RW)
0x1be: frame_vm_group_bin_12726 (RW)
0x1bf: frame_vm_group_bin_5656 (RW)
0x1c0: frame_vm_group_bin_21756 (RW)
0x1c1: frame_vm_group_bin_14582 (RW)
0x1c2: frame_vm_group_bin_7367 (RW)
0x1c3: frame_vm_group_bin_17499 (RW)
0x1c4: frame_vm_group_bin_16396 (RW)
0x1c5: frame_vm_group_bin_9215 (RW)
0x1c6: frame_vm_group_bin_2033 (RW)
0x1c7: frame_vm_group_bin_18129 (RW)
0x1c8: frame_vm_group_bin_11041 (RW)
0x1c9: frame_vm_group_bin_3856 (RW)
0x1c: frame_vm_group_bin_2800 (RW)
0x1ca: frame_vm_group_bin_19954 (RW)
0x1cb: frame_vm_group_bin_12753 (RW)
0x1cc: frame_vm_group_bin_5689 (RW)
0x1cd: frame_vm_group_bin_21788 (RW)
0x1ce: frame_vm_group_bin_14614 (RW)
0x1cf: frame_vm_group_bin_7400 (RW)
0x1d0: frame_vm_group_bin_22151 (RW)
0x1d1: frame_vm_group_bin_16429 (RW)
0x1d2: frame_vm_group_bin_9239 (RW)
0x1d3: frame_vm_group_bin_2066 (RW)
0x1d4: frame_vm_group_bin_18162 (RW)
0x1d5: frame_vm_group_bin_11074 (RW)
0x1d6: frame_vm_group_bin_3889 (RW)
0x1d7: frame_vm_group_bin_19987 (RW)
0x1d8: frame_vm_group_bin_12786 (RW)
0x1d9: frame_vm_group_bin_5722 (RW)
0x1d: frame_vm_group_bin_18874 (RW)
0x1da: frame_vm_group_bin_21823 (RW)
0x1db: frame_vm_group_bin_14648 (RW)
0x1dc: frame_vm_group_bin_7434 (RW)
0x1dd: frame_vm_group_bin_0283 (RW)
0x1de: frame_vm_group_bin_16463 (RW)
0x1df: frame_vm_group_bin_9263 (RW)
0x1e0: frame_vm_group_bin_2100 (RW)
0x1e1: frame_vm_group_bin_18195 (RW)
0x1e2: frame_vm_group_bin_11108 (RW)
0x1e3: frame_vm_group_bin_3923 (RW)
0x1e4: frame_vm_group_bin_20019 (RW)
0x1e5: frame_vm_group_bin_12819 (RW)
0x1e6: frame_vm_group_bin_5752 (RW)
0x1e7: frame_vm_group_bin_21856 (RW)
0x1e8: frame_vm_group_bin_14681 (RW)
0x1e9: frame_vm_group_bin_7467 (RW)
0x1e: frame_vm_group_bin_15178 (RW)
0x1ea: frame_vm_group_bin_0314 (RW)
0x1eb: frame_vm_group_bin_16496 (RW)
0x1ec: frame_vm_group_bin_9288 (RW)
0x1ed: frame_vm_group_bin_2134 (RW)
0x1ee: frame_vm_group_bin_18228 (RW)
0x1ef: frame_vm_group_bin_11140 (RW)
0x1f0: frame_vm_group_bin_3955 (RW)
0x1f1: frame_vm_group_bin_20052 (RW)
0x1f2: frame_vm_group_bin_12852 (RW)
0x1f3: frame_vm_group_bin_5775 (RW)
0x1f4: frame_vm_group_bin_21889 (RW)
0x1f5: frame_vm_group_bin_14714 (RW)
0x1f6: frame_vm_group_bin_7500 (RW)
0x1f7: frame_vm_group_bin_0345 (RW)
0x1f8: frame_vm_group_bin_16529 (RW)
0x1f9: frame_vm_group_bin_9317 (RW)
0x1f: frame_vm_group_bin_4612 (RW)
0x1fa: frame_vm_group_bin_2168 (RW)
0x1fb: frame_vm_group_bin_18262 (RW)
0x1fc: frame_vm_group_bin_11174 (RW)
0x1fd: frame_vm_group_bin_3989 (RW)
0x1fe: frame_vm_group_bin_20086 (RW)
0x1ff: frame_vm_group_bin_12886 (RW)
0x20: frame_vm_group_bin_20726 (RW)
0x21: frame_vm_group_bin_13527 (RW)
0x22: frame_vm_group_bin_6341 (RW)
0x23: frame_vm_group_bin_22534 (RW)
0x24: frame_vm_group_bin_15352 (RW)
0x25: frame_vm_group_bin_8161 (RW)
0x26: frame_vm_group_bin_1007 (RW)
0x27: frame_vm_group_bin_17198 (RW)
0x28: frame_vm_group_bin_9991 (RW)
0x29: frame_vm_group_bin_2833 (RW)
0x2: frame_vm_group_bin_2733 (RW)
0x2a: frame_vm_group_bin_18907 (RW)
0x2b: frame_vm_group_bin_19827 (RW)
0x2c: frame_vm_group_bin_4638 (RW)
0x2d: frame_vm_group_bin_20759 (RW)
0x2e: frame_vm_group_bin_13560 (RW)
0x2f: frame_vm_group_bin_6373 (RW)
0x30: frame_vm_group_bin_22567 (RW)
0x31: frame_vm_group_bin_15385 (RW)
0x32: frame_vm_group_bin_8194 (RW)
0x33: frame_vm_group_bin_1032 (RW)
0x34: frame_vm_group_bin_17231 (RW)
0x35: frame_vm_group_bin_10024 (RW)
0x36: frame_vm_group_bin_2865 (RW)
0x37: frame_vm_group_bin_18940 (RW)
0x38: frame_vm_group_bin_1177 (RW)
0x39: frame_vm_group_bin_4671 (RW)
0x3: frame_vm_group_bin_18806 (RW)
0x3a: frame_vm_group_bin_20793 (RW)
0x3b: frame_vm_group_bin_13594 (RW)
0x3c: frame_vm_group_bin_18730 (RW)
0x3d: frame_vm_group_bin_22601 (RW)
0x3e: frame_vm_group_bin_15419 (RW)
0x3f: frame_vm_group_bin_8228 (RW)
0x40: frame_vm_group_bin_1055 (RW)
0x41: frame_vm_group_bin_17264 (RW)
0x42: frame_vm_group_bin_10058 (RW)
0x43: frame_vm_group_bin_2901 (RW)
0x44: frame_vm_group_bin_18971 (RW)
0x45: frame_vm_group_bin_11830 (RW)
0x46: frame_vm_group_bin_4703 (RW)
0x47: frame_vm_group_bin_20825 (RW)
0x48: frame_vm_group_bin_13627 (RW)
0x49: frame_vm_group_bin_6437 (RW)
0x4: frame_vm_group_bin_11696 (RW)
0x4a: frame_vm_group_bin_22634 (RW)
0x4b: frame_vm_group_bin_15452 (RW)
0x4c: frame_vm_group_bin_8261 (RW)
0x4d: frame_vm_group_bin_1078 (RW)
0x4e: frame_vm_group_bin_17297 (RW)
0x4f: frame_vm_group_bin_10091 (RW)
0x50: frame_vm_group_bin_2934 (RW)
0x51: frame_vm_group_bin_19004 (RW)
0x52: frame_vm_group_bin_10561 (RW)
0x53: frame_vm_group_bin_4735 (RW)
0x54: frame_vm_group_bin_20854 (RW)
0x55: frame_vm_group_bin_13659 (RW)
0x56: frame_vm_group_bin_6470 (RW)
0x57: frame_vm_group_bin_22667 (RW)
0x58: frame_vm_group_bin_15485 (RW)
0x59: frame_vm_group_bin_8293 (RW)
0x5: frame_vm_group_bin_4563 (RW)
0x5a: frame_vm_group_bin_1106 (RW)
0x5b: frame_vm_group_bin_17331 (RW)
0x5c: frame_vm_group_bin_10125 (RW)
0x5d: frame_vm_group_bin_2968 (RW)
0x5e: frame_vm_group_bin_19038 (RW)
0x5f: frame_vm_group_bin_15202 (RW)
0x60: frame_vm_group_bin_4769 (RW)
0x61: frame_vm_group_bin_20880 (RW)
0x62: frame_vm_group_bin_13693 (RW)
0x63: frame_vm_group_bin_6504 (RW)
0x64: frame_vm_group_bin_22701 (RW)
0x65: frame_vm_group_bin_15518 (RW)
0x66: frame_vm_group_bin_8327 (RW)
0x67: frame_vm_group_bin_1138 (RW)
0x68: frame_vm_group_bin_17363 (RW)
0x69: frame_vm_group_bin_10160 (RW)
0x6: frame_vm_group_bin_20659 (RW)
0x6a: frame_vm_group_bin_3001 (RW)
0x6b: frame_vm_group_bin_19071 (RW)
0x6c: frame_vm_group_bin_19851 (RW)
0x6d: frame_vm_group_bin_4802 (RW)
0x6e: frame_vm_group_bin_20907 (RW)
0x6f: frame_vm_group_bin_13725 (RW)
0x70: frame_vm_group_bin_6537 (RW)
0x71: frame_vm_group_bin_22734 (RW)
0x72: frame_vm_group_bin_15550 (RW)
0x73: frame_vm_group_bin_8360 (RW)
0x74: frame_vm_group_bin_1171 (RW)
0x75: frame_vm_group_bin_17393 (RW)
0x76: frame_vm_group_bin_10193 (RW)
0x77: frame_vm_group_bin_3034 (RW)
0x78: frame_vm_group_bin_19104 (RW)
0x79: frame_vm_group_bin_1200 (RW)
0x7: frame_vm_group_bin_13460 (RW)
0x7a: frame_vm_group_bin_4835 (RW)
0x7b: frame_vm_group_bin_20936 (RW)
0x7c: frame_vm_group_bin_13760 (RW)
0x7d: frame_vm_group_bin_6571 (RW)
0x7e: frame_vm_group_bin_22767 (RW)
0x7f: frame_vm_group_bin_15584 (RW)
0x80: frame_vm_group_bin_8394 (RW)
0x81: frame_vm_group_bin_1205 (RW)
0x82: frame_vm_group_bin_17421 (RW)
0x83: frame_vm_group_bin_10227 (RW)
0x84: frame_vm_group_bin_3068 (RW)
0x85: frame_vm_group_bin_19136 (RW)
0x86: frame_vm_group_bin_11973 (RW)
0x87: frame_vm_group_bin_4868 (RW)
0x88: frame_vm_group_bin_20963 (RW)
0x89: frame_vm_group_bin_13793 (RW)
0x8: frame_vm_group_bin_6275 (RW)
0x8a: frame_vm_group_bin_6604 (RW)
0x8b: frame_vm_group_bin_22800 (RW)
0x8c: frame_vm_group_bin_15617 (RW)
0x8d: frame_vm_group_bin_8427 (RW)
0x8e: frame_vm_group_bin_1238 (RW)
0x8f: frame_vm_group_bin_17446 (RW)
0x90: frame_vm_group_bin_10260 (RW)
0x91: frame_vm_group_bin_3101 (RW)
0x92: frame_vm_group_bin_19169 (RW)
0x93: frame_vm_group_bin_12005 (RW)
0x94: frame_vm_group_bin_4901 (RW)
0x95: frame_vm_group_bin_20994 (RW)
0x96: frame_vm_group_bin_13824 (RW)
0x97: frame_vm_group_bin_6637 (RW)
0x98: frame_vm_group_bin_22833 (RW)
0x99: frame_vm_group_bin_15650 (RW)
0x9: frame_vm_group_bin_22468 (RW)
0x9a: frame_vm_group_bin_8461 (RW)
0x9b: frame_vm_group_bin_1271 (RW)
0x9c: frame_vm_group_bin_20952 (RW)
0x9d: frame_vm_group_bin_10294 (RW)
0x9e: frame_vm_group_bin_3134 (RW)
0x9f: frame_vm_group_bin_19203 (RW)
0xa0: frame_vm_group_bin_12036 (RW)
0xa1: frame_vm_group_bin_4933 (RW)
0xa2: frame_vm_group_bin_21028 (RW)
0xa3: frame_vm_group_bin_13855 (RW)
0xa4: frame_vm_group_bin_6671 (RW)
0xa5: frame_vm_group_bin_22867 (RW)
0xa6: frame_vm_group_bin_15684 (RW)
0xa7: frame_vm_group_bin_8494 (RW)
0xa8: frame_vm_group_bin_1302 (RW)
0xa9: frame_vm_group_bin_2324 (RW)
0xa: frame_vm_group_bin_15285 (RW)
0xaa: frame_vm_group_bin_10327 (RW)
0xab: frame_vm_group_bin_3167 (RW)
0xac: frame_vm_group_bin_19236 (RW)
0xad: frame_vm_group_bin_12063 (RW)
0xae: frame_vm_group_bin_4964 (RW)
0xaf: frame_vm_group_bin_21062 (RW)
0xb0: frame_vm_group_bin_13884 (RW)
0xb1: frame_vm_group_bin_6704 (RW)
0xb2: frame_vm_group_bin_22900 (RW)
0xb3: frame_vm_group_bin_15717 (RW)
0xb4: frame_vm_group_bin_8526 (RW)
0xb5: frame_vm_group_bin_1334 (RW)
0xb6: frame_vm_group_bin_6940 (RW)
0xb7: frame_vm_group_bin_10360 (RW)
0xb8: frame_vm_group_bin_3200 (RW)
0xb9: frame_vm_group_bin_19269 (RW)
0xb: frame_vm_group_bin_8095 (RW)
0xba: frame_vm_group_bin_12097 (RW)
0xbb: frame_vm_group_bin_4998 (RW)
0xbc: frame_vm_group_bin_21096 (RW)
0xbd: frame_vm_group_bin_13918 (RW)
0xbe: frame_vm_group_bin_6737 (RW)
0xbf: frame_vm_group_bin_22934 (RW)
0xc0: frame_vm_group_bin_15751 (RW)
0xc1: frame_vm_group_bin_8558 (RW)
0xc2: frame_vm_group_bin_1369 (RW)
0xc3: frame_vm_group_bin_11671 (RW)
0xc4: frame_vm_group_bin_10393 (RW)
0xc5: frame_vm_group_bin_3233 (RW)
0xc6: frame_vm_group_bin_19303 (RW)
0xc7: frame_vm_group_bin_12129 (RW)
0xc8: frame_vm_group_bin_5031 (RW)
0xc9: frame_vm_group_bin_21129 (RW)
0xc: frame_vm_group_bin_0940 (RW)
0xca: frame_vm_group_bin_13951 (RW)
0xcb: frame_vm_group_bin_6769 (RW)
0xcc: frame_vm_group_bin_22966 (RW)
0xcd: frame_vm_group_bin_15784 (RW)
0xce: frame_vm_group_bin_8591 (RW)
0xcf: frame_vm_group_bin_1402 (RW)
0xd0: frame_vm_group_bin_16342 (RW)
0xd1: frame_vm_group_bin_10418 (RW)
0xd2: frame_vm_group_bin_3266 (RW)
0xd3: frame_vm_group_bin_19336 (RW)
0xd4: frame_vm_group_bin_12161 (RW)
0xd5: frame_vm_group_bin_5064 (RW)
0xd6: frame_vm_group_bin_21161 (RW)
0xd7: frame_vm_group_bin_13984 (RW)
0xd8: frame_vm_group_bin_6802 (RW)
0xd9: frame_vm_group_bin_22999 (RW)
0xd: frame_vm_group_bin_17135 (RW)
0xda: frame_vm_group_bin_15817 (RW)
0xdb: frame_vm_group_bin_8624 (RW)
0xdc: frame_vm_group_bin_1436 (RW)
0xdd: frame_vm_group_bin_20975 (RW)
0xde: frame_vm_group_bin_10447 (RW)
0xdf: frame_vm_group_bin_3300 (RW)
0xe0: frame_vm_group_bin_19370 (RW)
0xe1: frame_vm_group_bin_12192 (RW)
0xe2: frame_vm_group_bin_5099 (RW)
0xe3: frame_vm_group_bin_21195 (RW)
0xe4: frame_vm_group_bin_14018 (RW)
0xe5: frame_vm_group_bin_6833 (RW)
0xe6: frame_vm_group_bin_23032 (RW)
0xe7: frame_vm_group_bin_15849 (RW)
0xe8: frame_vm_group_bin_8657 (RW)
0xe9: frame_vm_group_bin_1469 (RW)
0xe: frame_vm_group_bin_9926 (RW)
0xea: frame_vm_group_bin_2348 (RW)
0xeb: frame_vm_group_bin_10480 (RW)
0xec: frame_vm_group_bin_3333 (RW)
0xed: frame_vm_group_bin_19403 (RW)
0xee: frame_vm_group_bin_12222 (RW)
0xef: frame_vm_group_bin_5132 (RW)
0xf0: frame_vm_group_bin_21228 (RW)
0xf1: frame_vm_group_bin_14051 (RW)
0xf2: frame_vm_group_bin_6860 (RW)
0xf3: frame_vm_group_bin_23065 (RW)
0xf4: frame_vm_group_bin_15882 (RW)
0xf5: frame_vm_group_bin_8691 (RW)
0xf6: frame_vm_group_bin_1502 (RW)
0xf7: frame_vm_group_bin_17642 (RW)
0xf8: frame_vm_group_bin_10513 (RW)
0xf9: frame_vm_group_bin_3366 (RW)
0xf: frame_vm_group_bin_2766 (RW)
0xfa: frame_vm_group_bin_19436 (RW)
0xfb: frame_vm_group_bin_12255 (RW)
0xfc: frame_vm_group_bin_5166 (RW)
0xfd: frame_vm_group_bin_21262 (RW)
0xfe: frame_vm_group_bin_14085 (RW)
0xff: frame_vm_group_bin_6886 (RW)
}
pt_vm_group_bin_0115 {
0x0: frame_vm_group_bin_5074 (RW)
0x100: frame_vm_group_bin_11083 (RW)
0x101: frame_vm_group_bin_3898 (RW)
0x102: frame_vm_group_bin_19994 (RW)
0x103: frame_vm_group_bin_12795 (RW)
0x104: frame_vm_group_bin_5731 (RW)
0x105: frame_vm_group_bin_21831 (RW)
0x106: frame_vm_group_bin_14656 (RW)
0x107: frame_vm_group_bin_7442 (RW)
0x108: frame_vm_group_bin_0290 (RW)
0x109: frame_vm_group_bin_16471 (RW)
0x10: frame_vm_group_bin_6839 (RW)
0x10a: frame_vm_group_bin_9269 (RW)
0x10b: frame_vm_group_bin_2108 (RW)
0x10c: frame_vm_group_bin_18203 (RW)
0x10d: frame_vm_group_bin_11116 (RW)
0x10e: frame_vm_group_bin_3931 (RW)
0x10f: frame_vm_group_bin_20027 (RW)
0x110: frame_vm_group_bin_12827 (RW)
0x111: frame_vm_group_bin_5757 (RW)
0x112: frame_vm_group_bin_21864 (RW)
0x113: frame_vm_group_bin_14689 (RW)
0x114: frame_vm_group_bin_7475 (RW)
0x115: frame_vm_group_bin_0322 (RW)
0x116: frame_vm_group_bin_16504 (RW)
0x117: frame_vm_group_bin_9295 (RW)
0x118: frame_vm_group_bin_2142 (RW)
0x119: frame_vm_group_bin_18236 (RW)
0x11: frame_vm_group_bin_23040 (RW)
0x11a: frame_vm_group_bin_11149 (RW)
0x11b: frame_vm_group_bin_3964 (RW)
0x11c: frame_vm_group_bin_20061 (RW)
0x11d: frame_vm_group_bin_12861 (RW)
0x11e: frame_vm_group_bin_5782 (RW)
0x11f: frame_vm_group_bin_21898 (RW)
0x120: frame_vm_group_bin_14723 (RW)
0x121: frame_vm_group_bin_7508 (RW)
0x122: frame_vm_group_bin_0354 (RW)
0x123: frame_vm_group_bin_16538 (RW)
0x124: frame_vm_group_bin_9326 (RW)
0x125: frame_vm_group_bin_2176 (RW)
0x126: frame_vm_group_bin_18270 (RW)
0x127: frame_vm_group_bin_11182 (RW)
0x128: frame_vm_group_bin_3997 (RW)
0x129: frame_vm_group_bin_20094 (RW)
0x12: frame_vm_group_bin_15857 (RW)
0x12a: frame_vm_group_bin_12894 (RW)
0x12b: frame_vm_group_bin_14010 (RW)
0x12c: frame_vm_group_bin_21930 (RW)
0x12d: frame_vm_group_bin_14755 (RW)
0x12e: frame_vm_group_bin_7540 (RW)
0x12f: frame_vm_group_bin_0385 (RW)
0x130: frame_vm_group_bin_16570 (RW)
0x131: frame_vm_group_bin_9359 (RW)
0x132: frame_vm_group_bin_2207 (RW)
0x133: frame_vm_group_bin_18303 (RW)
0x134: frame_vm_group_bin_11215 (RW)
0x135: frame_vm_group_bin_4030 (RW)
0x136: frame_vm_group_bin_20126 (RW)
0x137: frame_vm_group_bin_12927 (RW)
0x138: frame_vm_group_bin_5824 (RW)
0x139: frame_vm_group_bin_21963 (RW)
0x13: frame_vm_group_bin_8665 (RW)
0x13a: frame_vm_group_bin_14788 (RW)
0x13b: frame_vm_group_bin_7573 (RW)
0x13c: frame_vm_group_bin_0415 (RW)
0x13d: frame_vm_group_bin_16603 (RW)
0x13e: frame_vm_group_bin_9394 (RW)
0x13f: frame_vm_group_bin_2236 (RW)
0x140: frame_vm_group_bin_18337 (RW)
0x141: frame_vm_group_bin_11249 (RW)
0x142: frame_vm_group_bin_4064 (RW)
0x143: frame_vm_group_bin_20159 (RW)
0x144: frame_vm_group_bin_12960 (RW)
0x145: frame_vm_group_bin_5849 (RW)
0x146: frame_vm_group_bin_21997 (RW)
0x147: frame_vm_group_bin_14821 (RW)
0x148: frame_vm_group_bin_7606 (RW)
0x149: frame_vm_group_bin_0446 (RW)
0x14: frame_vm_group_bin_1477 (RW)
0x14a: frame_vm_group_bin_16636 (RW)
0x14b: frame_vm_group_bin_9427 (RW)
0x14c: frame_vm_group_bin_2267 (RW)
0x14d: frame_vm_group_bin_18370 (RW)
0x14e: frame_vm_group_bin_11282 (RW)
0x14f: frame_vm_group_bin_4097 (RW)
0x150: frame_vm_group_bin_20191 (RW)
0x151: frame_vm_group_bin_12993 (RW)
0x152: frame_vm_group_bin_5875 (RW)
0x153: frame_vm_group_bin_22026 (RW)
0x154: frame_vm_group_bin_14854 (RW)
0x155: frame_vm_group_bin_7639 (RW)
0x156: frame_vm_group_bin_0479 (RW)
0x157: frame_vm_group_bin_16669 (RW)
0x158: frame_vm_group_bin_9460 (RW)
0x159: frame_vm_group_bin_2300 (RW)
0x15: frame_vm_group_bin_17617 (RW)
0x15a: frame_vm_group_bin_18403 (RW)
0x15b: frame_vm_group_bin_11316 (RW)
0x15c: frame_vm_group_bin_4130 (RW)
0x15d: frame_vm_group_bin_20225 (RW)
0x15e: frame_vm_group_bin_13029 (RW)
0x15f: frame_vm_group_bin_5902 (RW)
0x160: frame_vm_group_bin_22049 (RW)
0x161: frame_vm_group_bin_14888 (RW)
0x162: frame_vm_group_bin_7673 (RW)
0x163: frame_vm_group_bin_0512 (RW)
0x164: frame_vm_group_bin_16702 (RW)
0x165: frame_vm_group_bin_9494 (RW)
0x166: frame_vm_group_bin_2334 (RW)
0x167: frame_vm_group_bin_18435 (RW)
0x168: frame_vm_group_bin_11347 (RW)
0x169: frame_vm_group_bin_4162 (RW)
0x16: frame_vm_group_bin_10488 (RW)
0x16a: frame_vm_group_bin_20258 (RW)
0x16b: frame_vm_group_bin_13062 (RW)
0x16c: frame_vm_group_bin_14034 (RW)
0x16d: frame_vm_group_bin_22073 (RW)
0x16e: frame_vm_group_bin_14921 (RW)
0x16f: frame_vm_group_bin_7706 (RW)
0x170: frame_vm_group_bin_0544 (RW)
0x171: frame_vm_group_bin_16736 (RW)
0x172: frame_vm_group_bin_9527 (RW)
0x173: frame_vm_group_bin_2367 (RW)
0x174: frame_vm_group_bin_18466 (RW)
0x175: frame_vm_group_bin_11379 (RW)
0x176: frame_vm_group_bin_4195 (RW)
0x177: frame_vm_group_bin_20290 (RW)
0x178: frame_vm_group_bin_13095 (RW)
0x179: frame_vm_group_bin_18660 (RW)
0x17: frame_vm_group_bin_3341 (RW)
0x17a: frame_vm_group_bin_22104 (RW)
0x17b: frame_vm_group_bin_14955 (RW)
0x17c: frame_vm_group_bin_7739 (RW)
0x17d: frame_vm_group_bin_0576 (RW)
0x17e: frame_vm_group_bin_16770 (RW)
0x17f: frame_vm_group_bin_9561 (RW)
0x180: frame_vm_group_bin_2401 (RW)
0x181: frame_vm_group_bin_18495 (RW)
0x182: frame_vm_group_bin_11412 (RW)
0x183: frame_vm_group_bin_4228 (RW)
0x184: frame_vm_group_bin_20326 (RW)
0x185: frame_vm_group_bin_13129 (RW)
0x186: frame_vm_group_bin_5976 (RW)
0x187: frame_vm_group_bin_22137 (RW)
0x188: frame_vm_group_bin_14988 (RW)
0x189: frame_vm_group_bin_7772 (RW)
0x18: frame_vm_group_bin_19411 (RW)
0x18a: frame_vm_group_bin_0608 (RW)
0x18b: frame_vm_group_bin_16803 (RW)
0x18c: frame_vm_group_bin_9594 (RW)
0x18d: frame_vm_group_bin_2433 (RW)
0x18e: frame_vm_group_bin_18522 (RW)
0x18f: frame_vm_group_bin_11445 (RW)
0x190: frame_vm_group_bin_4261 (RW)
0x191: frame_vm_group_bin_20359 (RW)
0x192: frame_vm_group_bin_13162 (RW)
0x193: frame_vm_group_bin_6007 (RW)
0x194: frame_vm_group_bin_22170 (RW)
0x195: frame_vm_group_bin_15021 (RW)
0x196: frame_vm_group_bin_7805 (RW)
0x197: frame_vm_group_bin_0639 (RW)
0x198: frame_vm_group_bin_16836 (RW)
0x199: frame_vm_group_bin_9627 (RW)
0x19: frame_vm_group_bin_10724 (RW)
0x19a: frame_vm_group_bin_2467 (RW)
0x19b: frame_vm_group_bin_18547 (RW)
0x19c: frame_vm_group_bin_11479 (RW)
0x19d: frame_vm_group_bin_4295 (RW)
0x19e: frame_vm_group_bin_20393 (RW)
0x19f: frame_vm_group_bin_13196 (RW)
0x1: frame_vm_group_bin_21170 (RW)
0x1a0: frame_vm_group_bin_9391 (RW)
0x1a1: frame_vm_group_bin_22204 (RW)
0x1a2: frame_vm_group_bin_15050 (RW)
0x1a3: frame_vm_group_bin_7838 (RW)
0x1a4: frame_vm_group_bin_0674 (RW)
0x1a5: frame_vm_group_bin_16869 (RW)
0x1a6: frame_vm_group_bin_9661 (RW)
0x1a7: frame_vm_group_bin_2499 (RW)
0x1a8: frame_vm_group_bin_18576 (RW)
0x1a9: frame_vm_group_bin_11512 (RW)
0x1a: frame_vm_group_bin_5141 (RW)
0x1aa: frame_vm_group_bin_4328 (RW)
0x1ab: frame_vm_group_bin_20426 (RW)
0x1ac: frame_vm_group_bin_13229 (RW)
0x1ad: frame_vm_group_bin_14057 (RW)
0x1ae: frame_vm_group_bin_22237 (RW)
0x1af: frame_vm_group_bin_15074 (RW)
0x1b0: frame_vm_group_bin_7871 (RW)
0x1b1: frame_vm_group_bin_0707 (RW)
0x1b2: frame_vm_group_bin_16901 (RW)
0x1b3: frame_vm_group_bin_9693 (RW)
0x1b4: frame_vm_group_bin_2532 (RW)
0x1b5: frame_vm_group_bin_18609 (RW)
0x1b6: frame_vm_group_bin_11545 (RW)
0x1b7: frame_vm_group_bin_4363 (RW)
0x1b8: frame_vm_group_bin_20459 (RW)
0x1b9: frame_vm_group_bin_13262 (RW)
0x1b: frame_vm_group_bin_21237 (RW)
0x1ba: frame_vm_group_bin_6090 (RW)
0x1bb: frame_vm_group_bin_22271 (RW)
0x1bc: frame_vm_group_bin_15099 (RW)
0x1bd: frame_vm_group_bin_7905 (RW)
0x1be: frame_vm_group_bin_0741 (RW)
0x1bf: frame_vm_group_bin_16935 (RW)
0x1c0: frame_vm_group_bin_9727 (RW)
0x1c1: frame_vm_group_bin_2566 (RW)
0x1c2: frame_vm_group_bin_18642 (RW)
0x1c3: frame_vm_group_bin_11576 (RW)
0x1c4: frame_vm_group_bin_4397 (RW)
0x1c5: frame_vm_group_bin_20493 (RW)
0x1c6: frame_vm_group_bin_13296 (RW)
0x1c7: frame_vm_group_bin_6121 (RW)
0x1c8: frame_vm_group_bin_22303 (RW)
0x1c9: frame_vm_group_bin_15128 (RW)
0x1c: frame_vm_group_bin_14060 (RW)
0x1ca: frame_vm_group_bin_7939 (RW)
0x1cb: frame_vm_group_bin_0774 (RW)
0x1cc: frame_vm_group_bin_16968 (RW)
0x1cd: frame_vm_group_bin_9760 (RW)
0x1ce: frame_vm_group_bin_2599 (RW)
0x1cf: frame_vm_group_bin_18675 (RW)
0x1d0: frame_vm_group_bin_11601 (RW)
0x1d1: frame_vm_group_bin_4430 (RW)
0x1d2: frame_vm_group_bin_20526 (RW)
0x1d3: frame_vm_group_bin_13328 (RW)
0x1d4: frame_vm_group_bin_6153 (RW)
0x1d5: frame_vm_group_bin_22336 (RW)
0x1d6: frame_vm_group_bin_15151 (RW)
0x1d7: frame_vm_group_bin_7972 (RW)
0x1d8: frame_vm_group_bin_0807 (RW)
0x1d9: frame_vm_group_bin_17001 (RW)
0x1d: frame_vm_group_bin_6867 (RW)
0x1da: frame_vm_group_bin_9794 (RW)
0x1db: frame_vm_group_bin_2633 (RW)
0x1dc: frame_vm_group_bin_18708 (RW)
0x1dd: frame_vm_group_bin_21045 (RW)
0x1de: frame_vm_group_bin_4464 (RW)
0x1df: frame_vm_group_bin_20560 (RW)
0x1e0: frame_vm_group_bin_13362 (RW)
0x1e1: frame_vm_group_bin_6186 (RW)
0x1e2: frame_vm_group_bin_22369 (RW)
0x1e3: frame_vm_group_bin_15185 (RW)
0x1e4: frame_vm_group_bin_8004 (RW)
0x1e5: frame_vm_group_bin_0840 (RW)
0x1e6: frame_vm_group_bin_17035 (RW)
0x1e7: frame_vm_group_bin_9827 (RW)
0x1e8: frame_vm_group_bin_2666 (RW)
0x1e9: frame_vm_group_bin_18739 (RW)
0x1e: frame_vm_group_bin_23074 (RW)
0x1ea: frame_vm_group_bin_19804 (RW)
0x1eb: frame_vm_group_bin_4497 (RW)
0x1ec: frame_vm_group_bin_20593 (RW)
0x1ed: frame_vm_group_bin_13393 (RW)
0x1ee: frame_vm_group_bin_6213 (RW)
0x1ef: frame_vm_group_bin_22402 (RW)
0x1f0: frame_vm_group_bin_15218 (RW)
0x1f1: frame_vm_group_bin_8032 (RW)
0x1f2: frame_vm_group_bin_0873 (RW)
0x1f3: frame_vm_group_bin_17068 (RW)
0x1f4: frame_vm_group_bin_9860 (RW)
0x1f5: frame_vm_group_bin_2699 (RW)
0x1f6: frame_vm_group_bin_18772 (RW)
0x1f7: frame_vm_group_bin_1152 (RW)
0x1f8: frame_vm_group_bin_4530 (RW)
0x1f9: frame_vm_group_bin_20626 (RW)
0x1f: frame_vm_group_bin_15891 (RW)
0x1fa: frame_vm_group_bin_13427 (RW)
0x1fb: frame_vm_group_bin_18705 (RW)
0x1fc: frame_vm_group_bin_22435 (RW)
0x1fd: frame_vm_group_bin_15253 (RW)
0x1fe: frame_vm_group_bin_8063 (RW)
0x1ff: frame_vm_group_bin_0907 (RW)
0x20: frame_vm_group_bin_8700 (RW)
0x21: frame_vm_group_bin_1511 (RW)
0x22: frame_vm_group_bin_17651 (RW)
0x23: frame_vm_group_bin_10521 (RW)
0x24: frame_vm_group_bin_3374 (RW)
0x25: frame_vm_group_bin_19442 (RW)
0x26: frame_vm_group_bin_12263 (RW)
0x27: frame_vm_group_bin_5174 (RW)
0x28: frame_vm_group_bin_21270 (RW)
0x29: frame_vm_group_bin_14093 (RW)
0x2: frame_vm_group_bin_13993 (RW)
0x2a: frame_vm_group_bin_6892 (RW)
0x2b: frame_vm_group_bin_23107 (RW)
0x2c: frame_vm_group_bin_15924 (RW)
0x2d: frame_vm_group_bin_8733 (RW)
0x2e: frame_vm_group_bin_1544 (RW)
0x2f: frame_vm_group_bin_17682 (RW)
0x30: frame_vm_group_bin_10554 (RW)
0x31: frame_vm_group_bin_3403 (RW)
0x32: frame_vm_group_bin_19474 (RW)
0x33: frame_vm_group_bin_12296 (RW)
0x34: frame_vm_group_bin_5207 (RW)
0x35: frame_vm_group_bin_21303 (RW)
0x36: frame_vm_group_bin_14126 (RW)
0x37: frame_vm_group_bin_6916 (RW)
0x38: frame_vm_group_bin_23140 (RW)
0x39: frame_vm_group_bin_15957 (RW)
0x3: frame_vm_group_bin_6810 (RW)
0x3a: frame_vm_group_bin_8767 (RW)
0x3b: frame_vm_group_bin_1578 (RW)
0x3c: frame_vm_group_bin_7078 (RW)
0x3d: frame_vm_group_bin_10588 (RW)
0x3e: frame_vm_group_bin_3428 (RW)
0x3f: frame_vm_group_bin_19508 (RW)
0x40: frame_vm_group_bin_12329 (RW)
0x41: frame_vm_group_bin_5241 (RW)
0x42: frame_vm_group_bin_21335 (RW)
0x43: frame_vm_group_bin_14160 (RW)
0x44: frame_vm_group_bin_6947 (RW)
0x45: frame_vm_group_bin_23173 (RW)
0x46: frame_vm_group_bin_15993 (RW)
0x47: frame_vm_group_bin_8800 (RW)
0x48: frame_vm_group_bin_1611 (RW)
0x49: frame_vm_group_bin_11779 (RW)
0x4: frame_vm_group_bin_23007 (RW)
0x4a: frame_vm_group_bin_10621 (RW)
0x4b: frame_vm_group_bin_3450 (RW)
0x4c: frame_vm_group_bin_19541 (RW)
0x4d: frame_vm_group_bin_12362 (RW)
0x4e: frame_vm_group_bin_5274 (RW)
0x4f: frame_vm_group_bin_21368 (RW)
0x50: frame_vm_group_bin_14192 (RW)
0x51: frame_vm_group_bin_6979 (RW)
0x52: frame_vm_group_bin_23204 (RW)
0x53: frame_vm_group_bin_16026 (RW)
0x54: frame_vm_group_bin_8833 (RW)
0x55: frame_vm_group_bin_1644 (RW)
0x56: frame_vm_group_bin_17764 (RW)
0x57: frame_vm_group_bin_10653 (RW)
0x58: frame_vm_group_bin_3476 (RW)
0x59: frame_vm_group_bin_19575 (RW)
0x5: frame_vm_group_bin_15824 (RW)
0x5a: frame_vm_group_bin_12396 (RW)
0x5b: frame_vm_group_bin_5308 (RW)
0x5c: frame_vm_group_bin_21402 (RW)
0x5d: frame_vm_group_bin_14226 (RW)
0x5e: frame_vm_group_bin_7013 (RW)
0x5f: frame_vm_group_bin_23228 (RW)
0x60: frame_vm_group_bin_16060 (RW)
0x61: frame_vm_group_bin_8866 (RW)
0x62: frame_vm_group_bin_1678 (RW)
0x63: frame_vm_group_bin_17795 (RW)
0x64: frame_vm_group_bin_10686 (RW)
0x65: frame_vm_group_bin_3504 (RW)
0x66: frame_vm_group_bin_19609 (RW)
0x67: frame_vm_group_bin_12429 (RW)
0x68: frame_vm_group_bin_5339 (RW)
0x69: frame_vm_group_bin_21434 (RW)
0x6: frame_vm_group_bin_8632 (RW)
0x6a: frame_vm_group_bin_14258 (RW)
0x6b: frame_vm_group_bin_7045 (RW)
0x6c: frame_vm_group_bin_23249 (RW)
0x6d: frame_vm_group_bin_16092 (RW)
0x6e: frame_vm_group_bin_8898 (RW)
0x6f: frame_vm_group_bin_1710 (RW)
0x70: frame_vm_group_bin_17825 (RW)
0x71: frame_vm_group_bin_10718 (RW)
0x72: frame_vm_group_bin_3532 (RW)
0x73: frame_vm_group_bin_19640 (RW)
0x74: frame_vm_group_bin_12460 (RW)
0x75: frame_vm_group_bin_5370 (RW)
0x76: frame_vm_group_bin_21466 (RW)
0x77: frame_vm_group_bin_14290 (RW)
0x78: frame_vm_group_bin_7076 (RW)
0x79: frame_vm_group_bin_12834 (RW)
0x7: frame_vm_group_bin_1444 (RW)
0x7a: frame_vm_group_bin_16125 (RW)
0x7b: frame_vm_group_bin_8931 (RW)
0x7c: frame_vm_group_bin_1743 (RW)
0x7d: frame_vm_group_bin_7100 (RW)
0x7e: frame_vm_group_bin_10751 (RW)
0x7f: frame_vm_group_bin_3564 (RW)
0x80: frame_vm_group_bin_19668 (RW)
0x81: frame_vm_group_bin_12493 (RW)
0x82: frame_vm_group_bin_5403 (RW)
0x83: frame_vm_group_bin_21498 (RW)
0x84: frame_vm_group_bin_14322 (RW)
0x85: frame_vm_group_bin_7108 (RW)
0x86: frame_vm_group_bin_17551 (RW)
0x87: frame_vm_group_bin_16156 (RW)
0x88: frame_vm_group_bin_8963 (RW)
0x89: frame_vm_group_bin_1775 (RW)
0x8: frame_vm_group_bin_11762 (RW)
0x8a: frame_vm_group_bin_17879 (RW)
0x8b: frame_vm_group_bin_10783 (RW)
0x8c: frame_vm_group_bin_3598 (RW)
0x8d: frame_vm_group_bin_19698 (RW)
0x8e: frame_vm_group_bin_12526 (RW)
0x8f: frame_vm_group_bin_5436 (RW)
0x90: frame_vm_group_bin_21531 (RW)
0x91: frame_vm_group_bin_14355 (RW)
0x92: frame_vm_group_bin_7140 (RW)
0x93: frame_vm_group_bin_22223 (RW)
0x94: frame_vm_group_bin_16189 (RW)
0x95: frame_vm_group_bin_8996 (RW)
0x96: frame_vm_group_bin_1808 (RW)
0x97: frame_vm_group_bin_17910 (RW)
0x98: frame_vm_group_bin_10816 (RW)
0x99: frame_vm_group_bin_3631 (RW)
0x9: frame_vm_group_bin_10455 (RW)
0x9a: frame_vm_group_bin_19732 (RW)
0x9b: frame_vm_group_bin_12560 (RW)
0x9c: frame_vm_group_bin_5469 (RW)
0x9d: frame_vm_group_bin_21565 (RW)
0x9e: frame_vm_group_bin_14389 (RW)
0x9f: frame_vm_group_bin_7176 (RW)
0xa0: frame_vm_group_bin_0085 (RW)
0xa1: frame_vm_group_bin_16220 (RW)
0xa2: frame_vm_group_bin_9030 (RW)
0xa3: frame_vm_group_bin_1842 (RW)
0xa4: frame_vm_group_bin_17943 (RW)
0xa5: frame_vm_group_bin_10850 (RW)
0xa6: frame_vm_group_bin_3665 (RW)
0xa7: frame_vm_group_bin_19765 (RW)
0xa8: frame_vm_group_bin_12593 (RW)
0xa9: frame_vm_group_bin_5501 (RW)
0xa: frame_vm_group_bin_3308 (RW)
0xaa: frame_vm_group_bin_21598 (RW)
0xab: frame_vm_group_bin_14422 (RW)
0xac: frame_vm_group_bin_7209 (RW)
0xad: frame_vm_group_bin_8225 (RW)
0xae: frame_vm_group_bin_16246 (RW)
0xaf: frame_vm_group_bin_9063 (RW)
0xb0: frame_vm_group_bin_1875 (RW)
0xb1: frame_vm_group_bin_2513 (RW)
0xb2: frame_vm_group_bin_10882 (RW)
0xb3: frame_vm_group_bin_3698 (RW)
0xb4: frame_vm_group_bin_19798 (RW)
0xb5: frame_vm_group_bin_12626 (RW)
0xb6: frame_vm_group_bin_5533 (RW)
0xb7: frame_vm_group_bin_21631 (RW)
0xb8: frame_vm_group_bin_14455 (RW)
0xb9: frame_vm_group_bin_7242 (RW)
0xb: frame_vm_group_bin_19378 (RW)
0xba: frame_vm_group_bin_12858 (RW)
0xbb: frame_vm_group_bin_16274 (RW)
0xbc: frame_vm_group_bin_9097 (RW)
0xbd: frame_vm_group_bin_1909 (RW)
0xbe: frame_vm_group_bin_18007 (RW)
0xbf: frame_vm_group_bin_10917 (RW)
0xc0: frame_vm_group_bin_3732 (RW)
0xc1: frame_vm_group_bin_19832 (RW)
0xc2: frame_vm_group_bin_12658 (RW)
0xc3: frame_vm_group_bin_5567 (RW)
0xc4: frame_vm_group_bin_21665 (RW)
0xc5: frame_vm_group_bin_14489 (RW)
0xc6: frame_vm_group_bin_7276 (RW)
0xc7: frame_vm_group_bin_17567 (RW)
0xc8: frame_vm_group_bin_16305 (RW)
0xc9: frame_vm_group_bin_9130 (RW)
0xc: frame_vm_group_bin_12200 (RW)
0xca: frame_vm_group_bin_1942 (RW)
0xcb: frame_vm_group_bin_18040 (RW)
0xcc: frame_vm_group_bin_10950 (RW)
0xcd: frame_vm_group_bin_3765 (RW)
0xce: frame_vm_group_bin_19865 (RW)
0xcf: frame_vm_group_bin_12682 (RW)
0xd0: frame_vm_group_bin_5599 (RW)
0xd1: frame_vm_group_bin_21697 (RW)
0xd2: frame_vm_group_bin_14523 (RW)
0xd3: frame_vm_group_bin_7308 (RW)
0xd4: frame_vm_group_bin_0183 (RW)
0xd5: frame_vm_group_bin_16337 (RW)
0xd6: frame_vm_group_bin_9162 (RW)
0xd7: frame_vm_group_bin_1974 (RW)
0xd8: frame_vm_group_bin_18072 (RW)
0xd9: frame_vm_group_bin_10982 (RW)
0xd: frame_vm_group_bin_5107 (RW)
0xda: frame_vm_group_bin_3798 (RW)
0xdb: frame_vm_group_bin_19898 (RW)
0xdc: frame_vm_group_bin_12707 (RW)
0xdd: frame_vm_group_bin_5631 (RW)
0xde: frame_vm_group_bin_21731 (RW)
0xdf: frame_vm_group_bin_14557 (RW)
0xe0: frame_vm_group_bin_7342 (RW)
0xe1: frame_vm_group_bin_0215 (RW)
0xe2: frame_vm_group_bin_16371 (RW)
0xe3: frame_vm_group_bin_9194 (RW)
0xe4: frame_vm_group_bin_2008 (RW)
0xe5: frame_vm_group_bin_18104 (RW)
0xe6: frame_vm_group_bin_11016 (RW)
0xe7: frame_vm_group_bin_3831 (RW)
0xe8: frame_vm_group_bin_19929 (RW)
0xe9: frame_vm_group_bin_12733 (RW)
0xe: frame_vm_group_bin_21203 (RW)
0xea: frame_vm_group_bin_5664 (RW)
0xeb: frame_vm_group_bin_21764 (RW)
0xec: frame_vm_group_bin_14590 (RW)
0xed: frame_vm_group_bin_7375 (RW)
0xee: frame_vm_group_bin_8249 (RW)
0xef: frame_vm_group_bin_16404 (RW)
0xf0: frame_vm_group_bin_9221 (RW)
0xf1: frame_vm_group_bin_2041 (RW)
0xf2: frame_vm_group_bin_18137 (RW)
0xf3: frame_vm_group_bin_11049 (RW)
0xf4: frame_vm_group_bin_3864 (RW)
0xf5: frame_vm_group_bin_19962 (RW)
0xf6: frame_vm_group_bin_12761 (RW)
0xf7: frame_vm_group_bin_5697 (RW)
0xf8: frame_vm_group_bin_21796 (RW)
0xf9: frame_vm_group_bin_14622 (RW)
0xf: frame_vm_group_bin_14026 (RW)
0xfa: frame_vm_group_bin_7409 (RW)
0xfb: frame_vm_group_bin_0263 (RW)
0xfc: frame_vm_group_bin_16438 (RW)
0xfd: frame_vm_group_bin_9246 (RW)
0xfe: frame_vm_group_bin_2075 (RW)
0xff: frame_vm_group_bin_18171 (RW)
}
pt_vm_group_bin_0117 {
0x0: frame_vm_group_bin_7177 (RW)
0x100: frame_vm_group_bin_13197 (RW)
0x101: frame_vm_group_bin_6039 (RW)
0x102: frame_vm_group_bin_22205 (RW)
0x103: frame_vm_group_bin_15051 (RW)
0x104: frame_vm_group_bin_7839 (RW)
0x105: frame_vm_group_bin_0675 (RW)
0x106: frame_vm_group_bin_16870 (RW)
0x107: frame_vm_group_bin_9662 (RW)
0x108: frame_vm_group_bin_2500 (RW)
0x109: frame_vm_group_bin_18577 (RW)
0x10: frame_vm_group_bin_9064 (RW)
0x10a: frame_vm_group_bin_11513 (RW)
0x10b: frame_vm_group_bin_4329 (RW)
0x10c: frame_vm_group_bin_20427 (RW)
0x10d: frame_vm_group_bin_13230 (RW)
0x10e: frame_vm_group_bin_6062 (RW)
0x10f: frame_vm_group_bin_22238 (RW)
0x110: frame_vm_group_bin_6089 (RW)
0x111: frame_vm_group_bin_7872 (RW)
0x112: frame_vm_group_bin_0708 (RW)
0x113: frame_vm_group_bin_16902 (RW)
0x114: frame_vm_group_bin_9694 (RW)
0x115: frame_vm_group_bin_2533 (RW)
0x116: frame_vm_group_bin_18610 (RW)
0x117: frame_vm_group_bin_11546 (RW)
0x118: frame_vm_group_bin_4364 (RW)
0x119: frame_vm_group_bin_20460 (RW)
0x11: frame_vm_group_bin_1876 (RW)
0x11a: frame_vm_group_bin_13264 (RW)
0x11b: frame_vm_group_bin_6091 (RW)
0x11c: frame_vm_group_bin_12187 (RW)
0x11d: frame_vm_group_bin_15100 (RW)
0x11e: frame_vm_group_bin_7906 (RW)
0x11f: frame_vm_group_bin_0742 (RW)
0x120: frame_vm_group_bin_16936 (RW)
0x121: frame_vm_group_bin_9728 (RW)
0x122: frame_vm_group_bin_2567 (RW)
0x123: frame_vm_group_bin_18643 (RW)
0x124: frame_vm_group_bin_11577 (RW)
0x125: frame_vm_group_bin_4398 (RW)
0x126: frame_vm_group_bin_20494 (RW)
0x127: frame_vm_group_bin_13297 (RW)
0x128: frame_vm_group_bin_6122 (RW)
0x129: frame_vm_group_bin_22304 (RW)
0x12: frame_vm_group_bin_17974 (RW)
0x12a: frame_vm_group_bin_15464 (RW)
0x12b: frame_vm_group_bin_7940 (RW)
0x12c: frame_vm_group_bin_0775 (RW)
0x12d: frame_vm_group_bin_16969 (RW)
0x12e: frame_vm_group_bin_9761 (RW)
0x12f: frame_vm_group_bin_2600 (RW)
0x130: frame_vm_group_bin_18676 (RW)
0x131: frame_vm_group_bin_5466 (RW)
0x132: frame_vm_group_bin_4431 (RW)
0x133: frame_vm_group_bin_20527 (RW)
0x134: frame_vm_group_bin_13329 (RW)
0x135: frame_vm_group_bin_6154 (RW)
0x136: frame_vm_group_bin_22337 (RW)
0x137: frame_vm_group_bin_15152 (RW)
0x138: frame_vm_group_bin_7973 (RW)
0x139: frame_vm_group_bin_17306 (RW)
0x13: frame_vm_group_bin_10883 (RW)
0x13a: frame_vm_group_bin_17003 (RW)
0x13b: frame_vm_group_bin_9795 (RW)
0x13c: frame_vm_group_bin_2634 (RW)
0x13d: frame_vm_group_bin_18709 (RW)
0x13e: frame_vm_group_bin_14504 (RW)
0x13f: frame_vm_group_bin_4465 (RW)
0x140: frame_vm_group_bin_20561 (RW)
0x141: frame_vm_group_bin_13363 (RW)
0x142: frame_vm_group_bin_6187 (RW)
0x143: frame_vm_group_bin_22370 (RW)
0x144: frame_vm_group_bin_15186 (RW)
0x145: frame_vm_group_bin_8005 (RW)
0x146: frame_vm_group_bin_0841 (RW)
0x147: frame_vm_group_bin_17036 (RW)
0x148: frame_vm_group_bin_9828 (RW)
0x149: frame_vm_group_bin_2667 (RW)
0x14: frame_vm_group_bin_3699 (RW)
0x14a: frame_vm_group_bin_18740 (RW)
0x14b: frame_vm_group_bin_11649 (RW)
0x14c: frame_vm_group_bin_4498 (RW)
0x14d: frame_vm_group_bin_20594 (RW)
0x14e: frame_vm_group_bin_13394 (RW)
0x14f: frame_vm_group_bin_6214 (RW)
0x150: frame_vm_group_bin_22403 (RW)
0x151: frame_vm_group_bin_15219 (RW)
0x152: frame_vm_group_bin_4741 (RW)
0x153: frame_vm_group_bin_0874 (RW)
0x154: frame_vm_group_bin_17069 (RW)
0x155: frame_vm_group_bin_9861 (RW)
0x156: frame_vm_group_bin_2700 (RW)
0x157: frame_vm_group_bin_18773 (RW)
0x158: frame_vm_group_bin_11669 (RW)
0x159: frame_vm_group_bin_4531 (RW)
0x15: frame_vm_group_bin_19799 (RW)
0x15a: frame_vm_group_bin_20628 (RW)
0x15b: frame_vm_group_bin_13428 (RW)
0x15c: frame_vm_group_bin_6244 (RW)
0x15d: frame_vm_group_bin_22436 (RW)
0x15e: frame_vm_group_bin_15254 (RW)
0x15f: frame_vm_group_bin_8064 (RW)
0x160: frame_vm_group_bin_0908 (RW)
0x161: frame_vm_group_bin_17103 (RW)
0x162: frame_vm_group_bin_9894 (RW)
0x163: frame_vm_group_bin_2734 (RW)
0x164: frame_vm_group_bin_18807 (RW)
0x165: frame_vm_group_bin_11697 (RW)
0x166: frame_vm_group_bin_4564 (RW)
0x167: frame_vm_group_bin_20660 (RW)
0x168: frame_vm_group_bin_13461 (RW)
0x169: frame_vm_group_bin_6276 (RW)
0x16: frame_vm_group_bin_12627 (RW)
0x16a: frame_vm_group_bin_22469 (RW)
0x16b: frame_vm_group_bin_15286 (RW)
0x16c: frame_vm_group_bin_8096 (RW)
0x16d: frame_vm_group_bin_0941 (RW)
0x16e: frame_vm_group_bin_17136 (RW)
0x16f: frame_vm_group_bin_9927 (RW)
0x170: frame_vm_group_bin_2767 (RW)
0x171: frame_vm_group_bin_18841 (RW)
0x172: frame_vm_group_bin_11724 (RW)
0x173: frame_vm_group_bin_4035 (RW)
0x174: frame_vm_group_bin_20693 (RW)
0x175: frame_vm_group_bin_13494 (RW)
0x176: frame_vm_group_bin_6309 (RW)
0x177: frame_vm_group_bin_22502 (RW)
0x178: frame_vm_group_bin_15319 (RW)
0x179: frame_vm_group_bin_8128 (RW)
0x17: frame_vm_group_bin_5534 (RW)
0x17a: frame_vm_group_bin_0975 (RW)
0x17b: frame_vm_group_bin_17169 (RW)
0x17c: frame_vm_group_bin_9959 (RW)
0x17d: frame_vm_group_bin_2801 (RW)
0x17e: frame_vm_group_bin_18875 (RW)
0x17f: frame_vm_group_bin_11747 (RW)
0x180: frame_vm_group_bin_8673 (RW)
0x181: frame_vm_group_bin_20727 (RW)
0x182: frame_vm_group_bin_13528 (RW)
0x183: frame_vm_group_bin_6342 (RW)
0x184: frame_vm_group_bin_22535 (RW)
0x185: frame_vm_group_bin_15353 (RW)
0x186: frame_vm_group_bin_8162 (RW)
0x187: frame_vm_group_bin_1008 (RW)
0x188: frame_vm_group_bin_17199 (RW)
0x189: frame_vm_group_bin_9992 (RW)
0x18: frame_vm_group_bin_21632 (RW)
0x18a: frame_vm_group_bin_2834 (RW)
0x18b: frame_vm_group_bin_18908 (RW)
0x18c: frame_vm_group_bin_11770 (RW)
0x18d: frame_vm_group_bin_4639 (RW)
0x18e: frame_vm_group_bin_20760 (RW)
0x18f: frame_vm_group_bin_13561 (RW)
0x190: frame_vm_group_bin_6374 (RW)
0x191: frame_vm_group_bin_22568 (RW)
0x192: frame_vm_group_bin_15386 (RW)
0x193: frame_vm_group_bin_8195 (RW)
0x194: frame_vm_group_bin_1033 (RW)
0x195: frame_vm_group_bin_17232 (RW)
0x196: frame_vm_group_bin_10025 (RW)
0x197: frame_vm_group_bin_2866 (RW)
0x198: frame_vm_group_bin_18941 (RW)
0x199: frame_vm_group_bin_11797 (RW)
0x19: frame_vm_group_bin_14456 (RW)
0x19a: frame_vm_group_bin_4673 (RW)
0x19b: frame_vm_group_bin_20794 (RW)
0x19c: frame_vm_group_bin_13595 (RW)
0x19d: frame_vm_group_bin_6405 (RW)
0x19e: frame_vm_group_bin_22602 (RW)
0x19f: frame_vm_group_bin_15420 (RW)
0x1: frame_vm_group_bin_0086 (RW)
0x1a0: frame_vm_group_bin_8229 (RW)
0x1a1: frame_vm_group_bin_7952 (RW)
0x1a2: frame_vm_group_bin_17265 (RW)
0x1a3: frame_vm_group_bin_10059 (RW)
0x1a4: frame_vm_group_bin_2902 (RW)
0x1a5: frame_vm_group_bin_18972 (RW)
0x1a6: frame_vm_group_bin_11831 (RW)
0x1a7: frame_vm_group_bin_4704 (RW)
0x1a8: frame_vm_group_bin_20826 (RW)
0x1a9: frame_vm_group_bin_13628 (RW)
0x1a: frame_vm_group_bin_7244 (RW)
0x1aa: frame_vm_group_bin_6438 (RW)
0x1ab: frame_vm_group_bin_22635 (RW)
0x1ac: frame_vm_group_bin_15453 (RW)
0x1ad: frame_vm_group_bin_8262 (RW)
0x1ae: frame_vm_group_bin_12607 (RW)
0x1af: frame_vm_group_bin_17298 (RW)
0x1b0: frame_vm_group_bin_10092 (RW)
0x1b1: frame_vm_group_bin_2935 (RW)
0x1b2: frame_vm_group_bin_19005 (RW)
0x1b3: frame_vm_group_bin_11859 (RW)
0x1b4: frame_vm_group_bin_4736 (RW)
0x1b5: frame_vm_group_bin_20855 (RW)
0x1b6: frame_vm_group_bin_13660 (RW)
0x1b7: frame_vm_group_bin_6471 (RW)
0x1b8: frame_vm_group_bin_22668 (RW)
0x1b9: frame_vm_group_bin_15486 (RW)
0x1b: frame_vm_group_bin_0134 (RW)
0x1ba: frame_vm_group_bin_8295 (RW)
0x1bb: frame_vm_group_bin_1107 (RW)
0x1bc: frame_vm_group_bin_17332 (RW)
0x1bd: frame_vm_group_bin_10126 (RW)
0x1be: frame_vm_group_bin_2969 (RW)
0x1bf: frame_vm_group_bin_19039 (RW)
0x1c0: frame_vm_group_bin_11888 (RW)
0x1c1: frame_vm_group_bin_4770 (RW)
0x1c2: frame_vm_group_bin_7220 (RW)
0x1c3: frame_vm_group_bin_13694 (RW)
0x1c4: frame_vm_group_bin_6505 (RW)
0x1c5: frame_vm_group_bin_22702 (RW)
0x1c6: frame_vm_group_bin_15519 (RW)
0x1c7: frame_vm_group_bin_8328 (RW)
0x1c8: frame_vm_group_bin_1139 (RW)
0x1c9: frame_vm_group_bin_17364 (RW)
0x1c: frame_vm_group_bin_16275 (RW)
0x1ca: frame_vm_group_bin_10161 (RW)
0x1cb: frame_vm_group_bin_3002 (RW)
0x1cc: frame_vm_group_bin_19072 (RW)
0x1cd: frame_vm_group_bin_11911 (RW)
0x1ce: frame_vm_group_bin_4803 (RW)
0x1cf: frame_vm_group_bin_20908 (RW)
0x1d0: frame_vm_group_bin_13726 (RW)
0x1d1: frame_vm_group_bin_6538 (RW)
0x1d2: frame_vm_group_bin_22735 (RW)
0x1d3: frame_vm_group_bin_15551 (RW)
0x1d4: frame_vm_group_bin_8361 (RW)
0x1d5: frame_vm_group_bin_1172 (RW)
0x1d6: frame_vm_group_bin_17394 (RW)
0x1d7: frame_vm_group_bin_10194 (RW)
0x1d8: frame_vm_group_bin_3035 (RW)
0x1d9: frame_vm_group_bin_19105 (RW)
0x1d: frame_vm_group_bin_9098 (RW)
0x1da: frame_vm_group_bin_11941 (RW)
0x1db: frame_vm_group_bin_4836 (RW)
0x1dc: frame_vm_group_bin_20937 (RW)
0x1dd: frame_vm_group_bin_13761 (RW)
0x1de: frame_vm_group_bin_6572 (RW)
0x1df: frame_vm_group_bin_22768 (RW)
0x1e0: frame_vm_group_bin_15585 (RW)
0x1e1: frame_vm_group_bin_8395 (RW)
0x1e2: frame_vm_group_bin_1206 (RW)
0x1e3: frame_vm_group_bin_6521 (RW)
0x1e4: frame_vm_group_bin_10228 (RW)
0x1e5: frame_vm_group_bin_3069 (RW)
0x1e6: frame_vm_group_bin_19137 (RW)
0x1e7: frame_vm_group_bin_11974 (RW)
0x1e8: frame_vm_group_bin_4869 (RW)
0x1e9: frame_vm_group_bin_21259 (RW)
0x1e: frame_vm_group_bin_1910 (RW)
0x1ea: frame_vm_group_bin_13794 (RW)
0x1eb: frame_vm_group_bin_6605 (RW)
0x1ec: frame_vm_group_bin_22801 (RW)
0x1ed: frame_vm_group_bin_15618 (RW)
0x1ee: frame_vm_group_bin_8428 (RW)
0x1ef: frame_vm_group_bin_1239 (RW)
0x1f0: frame_vm_group_bin_11268 (RW)
0x1f1: frame_vm_group_bin_10261 (RW)
0x1f2: frame_vm_group_bin_3102 (RW)
0x1f3: frame_vm_group_bin_19170 (RW)
0x1f4: frame_vm_group_bin_12006 (RW)
0x1f5: frame_vm_group_bin_4902 (RW)
0x1f6: frame_vm_group_bin_20995 (RW)
0x1f7: frame_vm_group_bin_13825 (RW)
0x1f8: frame_vm_group_bin_6638 (RW)
0x1f9: frame_vm_group_bin_22834 (RW)
0x1f: frame_vm_group_bin_18008 (RW)
0x1fa: frame_vm_group_bin_15652 (RW)
0x1fb: frame_vm_group_bin_8462 (RW)
0x1fc: frame_vm_group_bin_17377 (RW)
0x1fd: frame_vm_group_bin_15911 (RW)
0x1fe: frame_vm_group_bin_10295 (RW)
0x1ff: frame_vm_group_bin_3135 (RW)
0x20: frame_vm_group_bin_10918 (RW)
0x21: frame_vm_group_bin_3733 (RW)
0x22: frame_vm_group_bin_19833 (RW)
0x23: frame_vm_group_bin_12659 (RW)
0x24: frame_vm_group_bin_5568 (RW)
0x25: frame_vm_group_bin_21666 (RW)
0x26: frame_vm_group_bin_14490 (RW)
0x27: frame_vm_group_bin_7277 (RW)
0x28: frame_vm_group_bin_0155 (RW)
0x29: frame_vm_group_bin_16306 (RW)
0x2: frame_vm_group_bin_16221 (RW)
0x2a: frame_vm_group_bin_9131 (RW)
0x2b: frame_vm_group_bin_1943 (RW)
0x2c: frame_vm_group_bin_18041 (RW)
0x2d: frame_vm_group_bin_10951 (RW)
0x2e: frame_vm_group_bin_3766 (RW)
0x2f: frame_vm_group_bin_19866 (RW)
0x30: frame_vm_group_bin_1018 (RW)
0x31: frame_vm_group_bin_5600 (RW)
0x32: frame_vm_group_bin_21698 (RW)
0x33: frame_vm_group_bin_14524 (RW)
0x34: frame_vm_group_bin_7309 (RW)
0x35: frame_vm_group_bin_0184 (RW)
0x36: frame_vm_group_bin_16338 (RW)
0x37: frame_vm_group_bin_9163 (RW)
0x38: frame_vm_group_bin_1975 (RW)
0x39: frame_vm_group_bin_18073 (RW)
0x3: frame_vm_group_bin_9031 (RW)
0x3a: frame_vm_group_bin_10984 (RW)
0x3b: frame_vm_group_bin_3799 (RW)
0x3c: frame_vm_group_bin_19899 (RW)
0x3d: frame_vm_group_bin_12708 (RW)
0x3e: frame_vm_group_bin_5632 (RW)
0x3f: frame_vm_group_bin_21732 (RW)
0x40: frame_vm_group_bin_14558 (RW)
0x41: frame_vm_group_bin_7343 (RW)
0x42: frame_vm_group_bin_0216 (RW)
0x43: frame_vm_group_bin_16372 (RW)
0x44: frame_vm_group_bin_9195 (RW)
0x45: frame_vm_group_bin_2009 (RW)
0x46: frame_vm_group_bin_18105 (RW)
0x47: frame_vm_group_bin_11017 (RW)
0x48: frame_vm_group_bin_3832 (RW)
0x49: frame_vm_group_bin_19930 (RW)
0x4: frame_vm_group_bin_1843 (RW)
0x4a: frame_vm_group_bin_10385 (RW)
0x4b: frame_vm_group_bin_5665 (RW)
0x4c: frame_vm_group_bin_21765 (RW)
0x4d: frame_vm_group_bin_14591 (RW)
0x4e: frame_vm_group_bin_7376 (RW)
0x4f: frame_vm_group_bin_0241 (RW)
0x50: frame_vm_group_bin_16405 (RW)
0x51: frame_vm_group_bin_0304 (RW)
0x52: frame_vm_group_bin_2042 (RW)
0x53: frame_vm_group_bin_18138 (RW)
0x54: frame_vm_group_bin_11050 (RW)
0x55: frame_vm_group_bin_3865 (RW)
0x56: frame_vm_group_bin_19963 (RW)
0x57: frame_vm_group_bin_12762 (RW)
0x58: frame_vm_group_bin_5698 (RW)
0x59: frame_vm_group_bin_21799 (RW)
0x5: frame_vm_group_bin_17944 (RW)
0x5a: frame_vm_group_bin_14624 (RW)
0x5b: frame_vm_group_bin_7410 (RW)
0x5c: frame_vm_group_bin_0264 (RW)
0x5d: frame_vm_group_bin_16439 (RW)
0x5e: frame_vm_group_bin_9247 (RW)
0x5f: frame_vm_group_bin_2076 (RW)
0x60: frame_vm_group_bin_18172 (RW)
0x61: frame_vm_group_bin_11084 (RW)
0x62: frame_vm_group_bin_3899 (RW)
0x63: frame_vm_group_bin_19995 (RW)
0x64: frame_vm_group_bin_12796 (RW)
0x65: frame_vm_group_bin_5732 (RW)
0x66: frame_vm_group_bin_21832 (RW)
0x67: frame_vm_group_bin_14657 (RW)
0x68: frame_vm_group_bin_7443 (RW)
0x69: frame_vm_group_bin_0291 (RW)
0x6: frame_vm_group_bin_10851 (RW)
0x6a: frame_vm_group_bin_16472 (RW)
0x6b: frame_vm_group_bin_9651 (RW)
0x6c: frame_vm_group_bin_2109 (RW)
0x6d: frame_vm_group_bin_18204 (RW)
0x6e: frame_vm_group_bin_11117 (RW)
0x6f: frame_vm_group_bin_3932 (RW)
0x70: frame_vm_group_bin_20028 (RW)
0x71: frame_vm_group_bin_12828 (RW)
0x72: frame_vm_group_bin_5758 (RW)
0x73: frame_vm_group_bin_21865 (RW)
0x74: frame_vm_group_bin_14690 (RW)
0x75: frame_vm_group_bin_7476 (RW)
0x76: frame_vm_group_bin_0323 (RW)
0x77: frame_vm_group_bin_16505 (RW)
0x78: frame_vm_group_bin_9296 (RW)
0x79: frame_vm_group_bin_2143 (RW)
0x7: frame_vm_group_bin_3666 (RW)
0x7a: frame_vm_group_bin_18238 (RW)
0x7b: frame_vm_group_bin_11150 (RW)
0x7c: frame_vm_group_bin_3965 (RW)
0x7d: frame_vm_group_bin_20062 (RW)
0x7e: frame_vm_group_bin_12862 (RW)
0x7f: frame_vm_group_bin_5783 (RW)
0x80: frame_vm_group_bin_21899 (RW)
0x81: frame_vm_group_bin_14724 (RW)
0x82: frame_vm_group_bin_7509 (RW)
0x83: frame_vm_group_bin_0355 (RW)
0x84: frame_vm_group_bin_16539 (RW)
0x85: frame_vm_group_bin_9327 (RW)
0x86: frame_vm_group_bin_2177 (RW)
0x87: frame_vm_group_bin_18271 (RW)
0x88: frame_vm_group_bin_11183 (RW)
0x89: frame_vm_group_bin_3998 (RW)
0x8: frame_vm_group_bin_19766 (RW)
0x8a: frame_vm_group_bin_20095 (RW)
0x8b: frame_vm_group_bin_12895 (RW)
0x8c: frame_vm_group_bin_5803 (RW)
0x8d: frame_vm_group_bin_21931 (RW)
0x8e: frame_vm_group_bin_14756 (RW)
0x8f: frame_vm_group_bin_7541 (RW)
0x90: frame_vm_group_bin_0386 (RW)
0x91: frame_vm_group_bin_16571 (RW)
0x92: frame_vm_group_bin_9360 (RW)
0x93: frame_vm_group_bin_2208 (RW)
0x94: frame_vm_group_bin_18304 (RW)
0x95: frame_vm_group_bin_11216 (RW)
0x96: frame_vm_group_bin_4031 (RW)
0x97: frame_vm_group_bin_20127 (RW)
0x98: frame_vm_group_bin_12928 (RW)
0x99: frame_vm_group_bin_5825 (RW)
0x9: frame_vm_group_bin_12594 (RW)
0x9a: frame_vm_group_bin_21965 (RW)
0x9b: frame_vm_group_bin_14789 (RW)
0x9c: frame_vm_group_bin_7574 (RW)
0x9d: frame_vm_group_bin_0416 (RW)
0x9e: frame_vm_group_bin_16604 (RW)
0x9f: frame_vm_group_bin_9395 (RW)
0xa0: frame_vm_group_bin_3586 (RW)
0xa1: frame_vm_group_bin_18338 (RW)
0xa2: frame_vm_group_bin_11250 (RW)
0xa3: frame_vm_group_bin_4065 (RW)
0xa4: frame_vm_group_bin_20160 (RW)
0xa5: frame_vm_group_bin_12961 (RW)
0xa6: frame_vm_group_bin_5850 (RW)
0xa7: frame_vm_group_bin_21998 (RW)
0xa8: frame_vm_group_bin_14822 (RW)
0xa9: frame_vm_group_bin_7607 (RW)
0xa: frame_vm_group_bin_5502 (RW)
0xaa: frame_vm_group_bin_0447 (RW)
0xab: frame_vm_group_bin_16637 (RW)
0xac: frame_vm_group_bin_9428 (RW)
0xad: frame_vm_group_bin_2268 (RW)
0xae: frame_vm_group_bin_18371 (RW)
0xaf: frame_vm_group_bin_11283 (RW)
0xb0: frame_vm_group_bin_4098 (RW)
0xb1: frame_vm_group_bin_20192 (RW)
0xb2: frame_vm_group_bin_12994 (RW)
0xb3: frame_vm_group_bin_5876 (RW)
0xb4: frame_vm_group_bin_22027 (RW)
0xb5: frame_vm_group_bin_14855 (RW)
0xb6: frame_vm_group_bin_7640 (RW)
0xb7: frame_vm_group_bin_0480 (RW)
0xb8: frame_vm_group_bin_16670 (RW)
0xb9: frame_vm_group_bin_9461 (RW)
0xb: frame_vm_group_bin_21599 (RW)
0xba: frame_vm_group_bin_2302 (RW)
0xbb: frame_vm_group_bin_18404 (RW)
0xbc: frame_vm_group_bin_11317 (RW)
0xbd: frame_vm_group_bin_4131 (RW)
0xbe: frame_vm_group_bin_20226 (RW)
0xbf: frame_vm_group_bin_13030 (RW)
0xc0: frame_vm_group_bin_5903 (RW)
0xc1: frame_vm_group_bin_2894 (RW)
0xc2: frame_vm_group_bin_14889 (RW)
0xc3: frame_vm_group_bin_7674 (RW)
0xc4: frame_vm_group_bin_0513 (RW)
0xc5: frame_vm_group_bin_16703 (RW)
0xc6: frame_vm_group_bin_9495 (RW)
0xc7: frame_vm_group_bin_2335 (RW)
0xc8: frame_vm_group_bin_18436 (RW)
0xc9: frame_vm_group_bin_11348 (RW)
0xc: frame_vm_group_bin_14423 (RW)
0xca: frame_vm_group_bin_4163 (RW)
0xcb: frame_vm_group_bin_20259 (RW)
0xcc: frame_vm_group_bin_13063 (RW)
0xcd: frame_vm_group_bin_5928 (RW)
0xce: frame_vm_group_bin_22074 (RW)
0xcf: frame_vm_group_bin_14922 (RW)
0xd0: frame_vm_group_bin_7707 (RW)
0xd1: frame_vm_group_bin_0545 (RW)
0xd2: frame_vm_group_bin_16737 (RW)
0xd3: frame_vm_group_bin_9528 (RW)
0xd4: frame_vm_group_bin_2368 (RW)
0xd5: frame_vm_group_bin_18467 (RW)
0xd6: frame_vm_group_bin_11380 (RW)
0xd7: frame_vm_group_bin_4196 (RW)
0xd8: frame_vm_group_bin_20291 (RW)
0xd9: frame_vm_group_bin_13096 (RW)
0xd: frame_vm_group_bin_7210 (RW)
0xda: frame_vm_group_bin_5950 (RW)
0xdb: frame_vm_group_bin_22105 (RW)
0xdc: frame_vm_group_bin_14956 (RW)
0xdd: frame_vm_group_bin_7740 (RW)
0xde: frame_vm_group_bin_0577 (RW)
0xdf: frame_vm_group_bin_16771 (RW)
0xe0: frame_vm_group_bin_9562 (RW)
0xe1: frame_vm_group_bin_2402 (RW)
0xe2: frame_vm_group_bin_2167 (RW)
0xe3: frame_vm_group_bin_11413 (RW)
0xe4: frame_vm_group_bin_4229 (RW)
0xe5: frame_vm_group_bin_20327 (RW)
0xe6: frame_vm_group_bin_13130 (RW)
0xe7: frame_vm_group_bin_5977 (RW)
0xe8: frame_vm_group_bin_22138 (RW)
0xe9: frame_vm_group_bin_14989 (RW)
0xe: frame_vm_group_bin_0111 (RW)
0xea: frame_vm_group_bin_7773 (RW)
0xeb: frame_vm_group_bin_0609 (RW)
0xec: frame_vm_group_bin_16804 (RW)
0xed: frame_vm_group_bin_9595 (RW)
0xee: frame_vm_group_bin_2434 (RW)
0xef: frame_vm_group_bin_6804 (RW)
0xf0: frame_vm_group_bin_11446 (RW)
0xf1: frame_vm_group_bin_4262 (RW)
0xf2: frame_vm_group_bin_20360 (RW)
0xf3: frame_vm_group_bin_13163 (RW)
0xf4: frame_vm_group_bin_6008 (RW)
0xf5: frame_vm_group_bin_22171 (RW)
0xf6: frame_vm_group_bin_15022 (RW)
0xf7: frame_vm_group_bin_7806 (RW)
0xf8: frame_vm_group_bin_0640 (RW)
0xf9: frame_vm_group_bin_16837 (RW)
0xf: frame_vm_group_bin_1718 (RW)
0xfa: frame_vm_group_bin_9629 (RW)
0xfb: frame_vm_group_bin_12883 (RW)
0xfc: frame_vm_group_bin_18548 (RW)
0xfd: frame_vm_group_bin_11480 (RW)
0xfe: frame_vm_group_bin_4296 (RW)
0xff: frame_vm_group_bin_20394 (RW)
}
pt_vm_group_bin_0123 {
0x0: frame_vm_group_bin_4347 (RW)
0x100: frame_vm_group_bin_10344 (RW)
0x101: frame_vm_group_bin_3184 (RW)
0x102: frame_vm_group_bin_19253 (RW)
0x103: frame_vm_group_bin_12080 (RW)
0x104: frame_vm_group_bin_4981 (RW)
0x105: frame_vm_group_bin_21079 (RW)
0x106: frame_vm_group_bin_13901 (RW)
0x107: frame_vm_group_bin_6720 (RW)
0x108: frame_vm_group_bin_22917 (RW)
0x109: frame_vm_group_bin_15734 (RW)
0x10: frame_vm_group_bin_6105 (RW)
0x10a: frame_vm_group_bin_8543 (RW)
0x10b: frame_vm_group_bin_1351 (RW)
0x10c: frame_vm_group_bin_17526 (RW)
0x10d: frame_vm_group_bin_10377 (RW)
0x10e: frame_vm_group_bin_3217 (RW)
0x10f: frame_vm_group_bin_19286 (RW)
0x110: frame_vm_group_bin_12112 (RW)
0x111: frame_vm_group_bin_5014 (RW)
0x112: frame_vm_group_bin_21112 (RW)
0x113: frame_vm_group_bin_13934 (RW)
0x114: frame_vm_group_bin_6753 (RW)
0x115: frame_vm_group_bin_22950 (RW)
0x116: frame_vm_group_bin_15767 (RW)
0x117: frame_vm_group_bin_8574 (RW)
0x118: frame_vm_group_bin_1385 (RW)
0x119: frame_vm_group_bin_17550 (RW)
0x11: frame_vm_group_bin_22286 (RW)
0x11a: frame_vm_group_bin_10405 (RW)
0x11b: frame_vm_group_bin_3250 (RW)
0x11c: frame_vm_group_bin_19320 (RW)
0x11d: frame_vm_group_bin_12146 (RW)
0x11e: frame_vm_group_bin_5048 (RW)
0x11f: frame_vm_group_bin_21145 (RW)
0x120: frame_vm_group_bin_13968 (RW)
0x121: frame_vm_group_bin_6786 (RW)
0x122: frame_vm_group_bin_22983 (RW)
0x123: frame_vm_group_bin_15800 (RW)
0x124: frame_vm_group_bin_8607 (RW)
0x125: frame_vm_group_bin_1419 (RW)
0x126: frame_vm_group_bin_21188 (RW)
0x127: frame_vm_group_bin_10433 (RW)
0x128: frame_vm_group_bin_3283 (RW)
0x129: frame_vm_group_bin_19353 (RW)
0x12: frame_vm_group_bin_15112 (RW)
0x12a: frame_vm_group_bin_12176 (RW)
0x12b: frame_vm_group_bin_5082 (RW)
0x12c: frame_vm_group_bin_21178 (RW)
0x12d: frame_vm_group_bin_14001 (RW)
0x12e: frame_vm_group_bin_6817 (RW)
0x12f: frame_vm_group_bin_23015 (RW)
0x130: frame_vm_group_bin_15832 (RW)
0x131: frame_vm_group_bin_8640 (RW)
0x132: frame_vm_group_bin_1452 (RW)
0x133: frame_vm_group_bin_2561 (RW)
0x134: frame_vm_group_bin_10463 (RW)
0x135: frame_vm_group_bin_3316 (RW)
0x136: frame_vm_group_bin_19386 (RW)
0x137: frame_vm_group_bin_12206 (RW)
0x138: frame_vm_group_bin_5115 (RW)
0x139: frame_vm_group_bin_21211 (RW)
0x13: frame_vm_group_bin_7921 (RW)
0x13a: frame_vm_group_bin_14035 (RW)
0x13b: frame_vm_group_bin_6846 (RW)
0x13c: frame_vm_group_bin_23049 (RW)
0x13d: frame_vm_group_bin_15866 (RW)
0x13e: frame_vm_group_bin_8676 (RW)
0x13f: frame_vm_group_bin_1486 (RW)
0x140: frame_vm_group_bin_17626 (RW)
0x141: frame_vm_group_bin_10497 (RW)
0x142: frame_vm_group_bin_3350 (RW)
0x143: frame_vm_group_bin_19419 (RW)
0x144: frame_vm_group_bin_12238 (RW)
0x145: frame_vm_group_bin_5149 (RW)
0x146: frame_vm_group_bin_21245 (RW)
0x147: frame_vm_group_bin_14068 (RW)
0x148: frame_vm_group_bin_6874 (RW)
0x149: frame_vm_group_bin_23082 (RW)
0x14: frame_vm_group_bin_0757 (RW)
0x14a: frame_vm_group_bin_15899 (RW)
0x14b: frame_vm_group_bin_8708 (RW)
0x14c: frame_vm_group_bin_1519 (RW)
0x14d: frame_vm_group_bin_17659 (RW)
0x14e: frame_vm_group_bin_10529 (RW)
0x14f: frame_vm_group_bin_3381 (RW)
0x150: frame_vm_group_bin_19450 (RW)
0x151: frame_vm_group_bin_12271 (RW)
0x152: frame_vm_group_bin_5182 (RW)
0x153: frame_vm_group_bin_21278 (RW)
0x154: frame_vm_group_bin_14101 (RW)
0x155: frame_vm_group_bin_6897 (RW)
0x156: frame_vm_group_bin_23115 (RW)
0x157: frame_vm_group_bin_15932 (RW)
0x158: frame_vm_group_bin_8741 (RW)
0x159: frame_vm_group_bin_1552 (RW)
0x15: frame_vm_group_bin_16951 (RW)
0x15a: frame_vm_group_bin_16577 (RW)
0x15b: frame_vm_group_bin_10563 (RW)
0x15c: frame_vm_group_bin_3409 (RW)
0x15d: frame_vm_group_bin_19483 (RW)
0x15e: frame_vm_group_bin_12305 (RW)
0x15f: frame_vm_group_bin_5216 (RW)
0x160: frame_vm_group_bin_21311 (RW)
0x161: frame_vm_group_bin_14135 (RW)
0x162: frame_vm_group_bin_6925 (RW)
0x163: frame_vm_group_bin_23148 (RW)
0x164: frame_vm_group_bin_15966 (RW)
0x165: frame_vm_group_bin_8775 (RW)
0x166: frame_vm_group_bin_1586 (RW)
0x167: frame_vm_group_bin_21212 (RW)
0x168: frame_vm_group_bin_10596 (RW)
0x169: frame_vm_group_bin_3434 (RW)
0x16: frame_vm_group_bin_9743 (RW)
0x16a: frame_vm_group_bin_19516 (RW)
0x16b: frame_vm_group_bin_12337 (RW)
0x16c: frame_vm_group_bin_5249 (RW)
0x16d: frame_vm_group_bin_21343 (RW)
0x16e: frame_vm_group_bin_14168 (RW)
0x16f: frame_vm_group_bin_6955 (RW)
0x170: frame_vm_group_bin_23181 (RW)
0x171: frame_vm_group_bin_16001 (RW)
0x172: frame_vm_group_bin_8808 (RW)
0x173: frame_vm_group_bin_1619 (RW)
0x174: frame_vm_group_bin_2585 (RW)
0x175: frame_vm_group_bin_10629 (RW)
0x176: frame_vm_group_bin_3456 (RW)
0x177: frame_vm_group_bin_19549 (RW)
0x178: frame_vm_group_bin_12370 (RW)
0x179: frame_vm_group_bin_5282 (RW)
0x17: frame_vm_group_bin_2582 (RW)
0x17a: frame_vm_group_bin_21377 (RW)
0x17b: frame_vm_group_bin_14201 (RW)
0x17c: frame_vm_group_bin_6988 (RW)
0x17d: frame_vm_group_bin_23211 (RW)
0x17e: frame_vm_group_bin_16035 (RW)
0x17f: frame_vm_group_bin_8842 (RW)
0x180: frame_vm_group_bin_1653 (RW)
0x181: frame_vm_group_bin_17772 (RW)
0x182: frame_vm_group_bin_10661 (RW)
0x183: frame_vm_group_bin_3485 (RW)
0x184: frame_vm_group_bin_19584 (RW)
0x185: frame_vm_group_bin_12404 (RW)
0x186: frame_vm_group_bin_5315 (RW)
0x187: frame_vm_group_bin_21410 (RW)
0x188: frame_vm_group_bin_14234 (RW)
0x189: frame_vm_group_bin_7021 (RW)
0x18: frame_vm_group_bin_18658 (RW)
0x18a: frame_vm_group_bin_23233 (RW)
0x18b: frame_vm_group_bin_16068 (RW)
0x18c: frame_vm_group_bin_8874 (RW)
0x18d: frame_vm_group_bin_1686 (RW)
0x18e: frame_vm_group_bin_17803 (RW)
0x18f: frame_vm_group_bin_10694 (RW)
0x190: frame_vm_group_bin_3511 (RW)
0x191: frame_vm_group_bin_19617 (RW)
0x192: frame_vm_group_bin_12436 (RW)
0x193: frame_vm_group_bin_5347 (RW)
0x194: frame_vm_group_bin_21442 (RW)
0x195: frame_vm_group_bin_14266 (RW)
0x196: frame_vm_group_bin_7053 (RW)
0x197: frame_vm_group_bin_23254 (RW)
0x198: frame_vm_group_bin_16100 (RW)
0x199: frame_vm_group_bin_8906 (RW)
0x19: frame_vm_group_bin_11587 (RW)
0x19a: frame_vm_group_bin_1719 (RW)
0x19b: frame_vm_group_bin_16600 (RW)
0x19c: frame_vm_group_bin_10727 (RW)
0x19d: frame_vm_group_bin_3541 (RW)
0x19e: frame_vm_group_bin_19649 (RW)
0x19f: frame_vm_group_bin_12469 (RW)
0x1: frame_vm_group_bin_20443 (RW)
0x1a0: frame_vm_group_bin_5379 (RW)
0x1a1: frame_vm_group_bin_21475 (RW)
0x1a2: frame_vm_group_bin_14298 (RW)
0x1a3: frame_vm_group_bin_7085 (RW)
0x1a4: frame_vm_group_bin_3679 (RW)
0x1a5: frame_vm_group_bin_16132 (RW)
0x1a6: frame_vm_group_bin_8939 (RW)
0x1a7: frame_vm_group_bin_1751 (RW)
0x1a8: frame_vm_group_bin_21235 (RW)
0x1a9: frame_vm_group_bin_10759 (RW)
0x1a: frame_vm_group_bin_4414 (RW)
0x1aa: frame_vm_group_bin_3572 (RW)
0x1ab: frame_vm_group_bin_19676 (RW)
0x1ac: frame_vm_group_bin_12501 (RW)
0x1ad: frame_vm_group_bin_5411 (RW)
0x1ae: frame_vm_group_bin_21506 (RW)
0x1af: frame_vm_group_bin_14330 (RW)
0x1b0: frame_vm_group_bin_7116 (RW)
0x1b1: frame_vm_group_bin_8317 (RW)
0x1b2: frame_vm_group_bin_16164 (RW)
0x1b3: frame_vm_group_bin_8971 (RW)
0x1b4: frame_vm_group_bin_1783 (RW)
0x1b5: frame_vm_group_bin_17887 (RW)
0x1b6: frame_vm_group_bin_10791 (RW)
0x1b7: frame_vm_group_bin_3606 (RW)
0x1b8: frame_vm_group_bin_19706 (RW)
0x1b9: frame_vm_group_bin_12534 (RW)
0x1b: frame_vm_group_bin_20510 (RW)
0x1ba: frame_vm_group_bin_5445 (RW)
0x1bb: frame_vm_group_bin_21540 (RW)
0x1bc: frame_vm_group_bin_14364 (RW)
0x1bd: frame_vm_group_bin_7149 (RW)
0x1be: frame_vm_group_bin_12952 (RW)
0x1bf: frame_vm_group_bin_16198 (RW)
0x1c0: frame_vm_group_bin_9005 (RW)
0x1c1: frame_vm_group_bin_1817 (RW)
0x1c2: frame_vm_group_bin_17919 (RW)
0x1c3: frame_vm_group_bin_10825 (RW)
0x1c4: frame_vm_group_bin_3640 (RW)
0x1c5: frame_vm_group_bin_19740 (RW)
0x1c6: frame_vm_group_bin_12568 (RW)
0x1c7: frame_vm_group_bin_5476 (RW)
0x1c8: frame_vm_group_bin_21573 (RW)
0x1c9: frame_vm_group_bin_14397 (RW)
0x1c: frame_vm_group_bin_13313 (RW)
0x1ca: frame_vm_group_bin_7184 (RW)
0x1cb: frame_vm_group_bin_0091 (RW)
0x1cc: frame_vm_group_bin_16225 (RW)
0x1cd: frame_vm_group_bin_9038 (RW)
0x1ce: frame_vm_group_bin_1850 (RW)
0x1cf: frame_vm_group_bin_17950 (RW)
0x1d0: frame_vm_group_bin_10858 (RW)
0x1d1: frame_vm_group_bin_3673 (RW)
0x1d2: frame_vm_group_bin_19773 (RW)
0x1d3: frame_vm_group_bin_12601 (RW)
0x1d4: frame_vm_group_bin_5509 (RW)
0x1d5: frame_vm_group_bin_21606 (RW)
0x1d6: frame_vm_group_bin_14430 (RW)
0x1d7: frame_vm_group_bin_7217 (RW)
0x1d8: frame_vm_group_bin_0116 (RW)
0x1d9: frame_vm_group_bin_16251 (RW)
0x1d: frame_vm_group_bin_6138 (RW)
0x1da: frame_vm_group_bin_9072 (RW)
0x1db: frame_vm_group_bin_1884 (RW)
0x1dc: frame_vm_group_bin_17982 (RW)
0x1dd: frame_vm_group_bin_10892 (RW)
0x1de: frame_vm_group_bin_3707 (RW)
0x1df: frame_vm_group_bin_19807 (RW)
0x1e0: frame_vm_group_bin_12635 (RW)
0x1e1: frame_vm_group_bin_5542 (RW)
0x1e2: frame_vm_group_bin_21640 (RW)
0x1e3: frame_vm_group_bin_14464 (RW)
0x1e4: frame_vm_group_bin_7251 (RW)
0x1e5: frame_vm_group_bin_3704 (RW)
0x1e6: frame_vm_group_bin_16282 (RW)
0x1e7: frame_vm_group_bin_9105 (RW)
0x1e8: frame_vm_group_bin_1917 (RW)
0x1e9: frame_vm_group_bin_18015 (RW)
0x1e: frame_vm_group_bin_22320 (RW)
0x1ea: frame_vm_group_bin_10925 (RW)
0x1eb: frame_vm_group_bin_3740 (RW)
0x1ec: frame_vm_group_bin_19840 (RW)
0x1ed: frame_vm_group_bin_12664 (RW)
0x1ee: frame_vm_group_bin_5575 (RW)
0x1ef: frame_vm_group_bin_21673 (RW)
0x1f0: frame_vm_group_bin_14497 (RW)
0x1f1: frame_vm_group_bin_7284 (RW)
0x1f2: frame_vm_group_bin_8341 (RW)
0x1f3: frame_vm_group_bin_16313 (RW)
0x1f4: frame_vm_group_bin_9138 (RW)
0x1f5: frame_vm_group_bin_1950 (RW)
0x1f6: frame_vm_group_bin_18048 (RW)
0x1f7: frame_vm_group_bin_10958 (RW)
0x1f8: frame_vm_group_bin_3773 (RW)
0x1f9: frame_vm_group_bin_19873 (RW)
0x1f: frame_vm_group_bin_15139 (RW)
0x1fa: frame_vm_group_bin_12688 (RW)
0x1fb: frame_vm_group_bin_5608 (RW)
0x1fc: frame_vm_group_bin_21706 (RW)
0x1fd: frame_vm_group_bin_14532 (RW)
0x1fe: frame_vm_group_bin_7317 (RW)
0x1ff: frame_vm_group_bin_12976 (RW)
0x20: frame_vm_group_bin_7956 (RW)
0x21: frame_vm_group_bin_0791 (RW)
0x22: frame_vm_group_bin_16985 (RW)
0x23: frame_vm_group_bin_9777 (RW)
0x24: frame_vm_group_bin_2616 (RW)
0x25: frame_vm_group_bin_18692 (RW)
0x26: frame_vm_group_bin_11615 (RW)
0x27: frame_vm_group_bin_4447 (RW)
0x28: frame_vm_group_bin_20543 (RW)
0x29: frame_vm_group_bin_13345 (RW)
0x2: frame_vm_group_bin_13246 (RW)
0x2a: frame_vm_group_bin_6170 (RW)
0x2b: frame_vm_group_bin_22352 (RW)
0x2c: frame_vm_group_bin_15168 (RW)
0x2d: frame_vm_group_bin_7988 (RW)
0x2e: frame_vm_group_bin_0823 (RW)
0x2f: frame_vm_group_bin_17018 (RW)
0x30: frame_vm_group_bin_9810 (RW)
0x31: frame_vm_group_bin_2649 (RW)
0x32: frame_vm_group_bin_18724 (RW)
0x33: frame_vm_group_bin_20012 (RW)
0x34: frame_vm_group_bin_4480 (RW)
0x35: frame_vm_group_bin_20576 (RW)
0x36: frame_vm_group_bin_13377 (RW)
0x37: frame_vm_group_bin_6201 (RW)
0x38: frame_vm_group_bin_22385 (RW)
0x39: frame_vm_group_bin_15201 (RW)
0x3: frame_vm_group_bin_18896 (RW)
0x3a: frame_vm_group_bin_8019 (RW)
0x3b: frame_vm_group_bin_0857 (RW)
0x3c: frame_vm_group_bin_17052 (RW)
0x3d: frame_vm_group_bin_9844 (RW)
0x3e: frame_vm_group_bin_2683 (RW)
0x3f: frame_vm_group_bin_18756 (RW)
0x40: frame_vm_group_bin_1364 (RW)
0x41: frame_vm_group_bin_4514 (RW)
0x42: frame_vm_group_bin_20610 (RW)
0x43: frame_vm_group_bin_13410 (RW)
0x44: frame_vm_group_bin_6228 (RW)
0x45: frame_vm_group_bin_22418 (RW)
0x46: frame_vm_group_bin_15236 (RW)
0x47: frame_vm_group_bin_8048 (RW)
0x48: frame_vm_group_bin_0890 (RW)
0x49: frame_vm_group_bin_17085 (RW)
0x4: frame_vm_group_bin_22254 (RW)
0x4a: frame_vm_group_bin_9877 (RW)
0x4b: frame_vm_group_bin_2716 (RW)
0x4c: frame_vm_group_bin_18789 (RW)
0x4d: frame_vm_group_bin_11682 (RW)
0x4e: frame_vm_group_bin_4547 (RW)
0x4f: frame_vm_group_bin_20643 (RW)
0x50: frame_vm_group_bin_13443 (RW)
0x51: frame_vm_group_bin_6259 (RW)
0x52: frame_vm_group_bin_22451 (RW)
0x53: frame_vm_group_bin_15269 (RW)
0x54: frame_vm_group_bin_8079 (RW)
0x55: frame_vm_group_bin_0923 (RW)
0x56: frame_vm_group_bin_17118 (RW)
0x57: frame_vm_group_bin_9909 (RW)
0x58: frame_vm_group_bin_2749 (RW)
0x59: frame_vm_group_bin_18824 (RW)
0x5: frame_vm_group_bin_15088 (RW)
0x5a: frame_vm_group_bin_10748 (RW)
0x5b: frame_vm_group_bin_4576 (RW)
0x5c: frame_vm_group_bin_20676 (RW)
0x5d: frame_vm_group_bin_13477 (RW)
0x5e: frame_vm_group_bin_6292 (RW)
0x5f: frame_vm_group_bin_22485 (RW)
0x60: frame_vm_group_bin_15302 (RW)
0x61: frame_vm_group_bin_8111 (RW)
0x62: frame_vm_group_bin_0957 (RW)
0x63: frame_vm_group_bin_17151 (RW)
0x64: frame_vm_group_bin_9941 (RW)
0x65: frame_vm_group_bin_2783 (RW)
0x66: frame_vm_group_bin_18857 (RW)
0x67: frame_vm_group_bin_15391 (RW)
0x68: frame_vm_group_bin_4600 (RW)
0x69: frame_vm_group_bin_20709 (RW)
0x6: frame_vm_group_bin_7888 (RW)
0x6a: frame_vm_group_bin_13510 (RW)
0x6b: frame_vm_group_bin_6324 (RW)
0x6c: frame_vm_group_bin_22518 (RW)
0x6d: frame_vm_group_bin_15335 (RW)
0x6e: frame_vm_group_bin_8144 (RW)
0x6f: frame_vm_group_bin_0990 (RW)
0x70: frame_vm_group_bin_17183 (RW)
0x71: frame_vm_group_bin_9974 (RW)
0x72: frame_vm_group_bin_2816 (RW)
0x73: frame_vm_group_bin_18890 (RW)
0x74: frame_vm_group_bin_20035 (RW)
0x75: frame_vm_group_bin_4624 (RW)
0x76: frame_vm_group_bin_20742 (RW)
0x77: frame_vm_group_bin_13543 (RW)
0x78: frame_vm_group_bin_6357 (RW)
0x79: frame_vm_group_bin_22550 (RW)
0x7: frame_vm_group_bin_0724 (RW)
0x7a: frame_vm_group_bin_15369 (RW)
0x7b: frame_vm_group_bin_8178 (RW)
0x7c: frame_vm_group_bin_1021 (RW)
0x7d: frame_vm_group_bin_17215 (RW)
0x7e: frame_vm_group_bin_10008 (RW)
0x7f: frame_vm_group_bin_2850 (RW)
0x80: frame_vm_group_bin_18924 (RW)
0x81: frame_vm_group_bin_11782 (RW)
0x82: frame_vm_group_bin_4655 (RW)
0x83: frame_vm_group_bin_20776 (RW)
0x84: frame_vm_group_bin_13577 (RW)
0x85: frame_vm_group_bin_6388 (RW)
0x86: frame_vm_group_bin_22584 (RW)
0x87: frame_vm_group_bin_15402 (RW)
0x88: frame_vm_group_bin_8211 (RW)
0x89: frame_vm_group_bin_1044 (RW)
0x8: frame_vm_group_bin_16918 (RW)
0x8a: frame_vm_group_bin_17247 (RW)
0x8b: frame_vm_group_bin_10041 (RW)
0x8c: frame_vm_group_bin_2884 (RW)
0x8d: frame_vm_group_bin_18956 (RW)
0x8e: frame_vm_group_bin_11813 (RW)
0x8f: frame_vm_group_bin_4687 (RW)
0x90: frame_vm_group_bin_20809 (RW)
0x91: frame_vm_group_bin_13610 (RW)
0x92: frame_vm_group_bin_6420 (RW)
0x93: frame_vm_group_bin_22617 (RW)
0x94: frame_vm_group_bin_15435 (RW)
0x95: frame_vm_group_bin_8244 (RW)
0x96: frame_vm_group_bin_1065 (RW)
0x97: frame_vm_group_bin_17280 (RW)
0x98: frame_vm_group_bin_10074 (RW)
0x99: frame_vm_group_bin_2917 (RW)
0x9: frame_vm_group_bin_9710 (RW)
0x9a: frame_vm_group_bin_18988 (RW)
0x9b: frame_vm_group_bin_11844 (RW)
0x9c: frame_vm_group_bin_4720 (RW)
0x9d: frame_vm_group_bin_20842 (RW)
0x9e: frame_vm_group_bin_13643 (RW)
0x9f: frame_vm_group_bin_5045 (RW)
0xa0: frame_vm_group_bin_22651 (RW)
0xa1: frame_vm_group_bin_15469 (RW)
0xa2: frame_vm_group_bin_8277 (RW)
0xa3: frame_vm_group_bin_1093 (RW)
0xa4: frame_vm_group_bin_17314 (RW)
0xa5: frame_vm_group_bin_10108 (RW)
0xa6: frame_vm_group_bin_2951 (RW)
0xa7: frame_vm_group_bin_19021 (RW)
0xa8: frame_vm_group_bin_15416 (RW)
0xa9: frame_vm_group_bin_4752 (RW)
0xa: frame_vm_group_bin_2549 (RW)
0xaa: frame_vm_group_bin_20867 (RW)
0xab: frame_vm_group_bin_13676 (RW)
0xac: frame_vm_group_bin_6487 (RW)
0xad: frame_vm_group_bin_22684 (RW)
0xae: frame_vm_group_bin_15502 (RW)
0xaf: frame_vm_group_bin_8310 (RW)
0xb0: frame_vm_group_bin_1121 (RW)
0xb1: frame_vm_group_bin_17347 (RW)
0xb2: frame_vm_group_bin_10141 (RW)
0xb3: frame_vm_group_bin_2984 (RW)
0xb4: frame_vm_group_bin_19054 (RW)
0xb5: frame_vm_group_bin_20058 (RW)
0xb6: frame_vm_group_bin_4785 (RW)
0xb7: frame_vm_group_bin_20893 (RW)
0xb8: frame_vm_group_bin_13709 (RW)
0xb9: frame_vm_group_bin_6520 (RW)
0xb: frame_vm_group_bin_18626 (RW)
0xba: frame_vm_group_bin_22718 (RW)
0xbb: frame_vm_group_bin_15535 (RW)
0xbc: frame_vm_group_bin_8344 (RW)
0xbd: frame_vm_group_bin_1155 (RW)
0xbe: frame_vm_group_bin_17380 (RW)
0xbf: frame_vm_group_bin_10177 (RW)
0xc0: frame_vm_group_bin_3018 (RW)
0xc1: frame_vm_group_bin_19088 (RW)
0xc2: frame_vm_group_bin_11926 (RW)
0xc3: frame_vm_group_bin_4818 (RW)
0xc4: frame_vm_group_bin_20922 (RW)
0xc5: frame_vm_group_bin_13742 (RW)
0xc6: frame_vm_group_bin_6554 (RW)
0xc7: frame_vm_group_bin_22750 (RW)
0xc8: frame_vm_group_bin_15567 (RW)
0xc9: frame_vm_group_bin_8377 (RW)
0xc: frame_vm_group_bin_11560 (RW)
0xca: frame_vm_group_bin_1188 (RW)
0xcb: frame_vm_group_bin_17408 (RW)
0xcc: frame_vm_group_bin_10210 (RW)
0xcd: frame_vm_group_bin_3051 (RW)
0xce: frame_vm_group_bin_19120 (RW)
0xcf: frame_vm_group_bin_11956 (RW)
0xd0: frame_vm_group_bin_4851 (RW)
0xd1: frame_vm_group_bin_20949 (RW)
0xd2: frame_vm_group_bin_13776 (RW)
0xd3: frame_vm_group_bin_6587 (RW)
0xd4: frame_vm_group_bin_22783 (RW)
0xd5: frame_vm_group_bin_15600 (RW)
0xd6: frame_vm_group_bin_8410 (RW)
0xd7: frame_vm_group_bin_1221 (RW)
0xd8: frame_vm_group_bin_17432 (RW)
0xd9: frame_vm_group_bin_10243 (RW)
0xd: frame_vm_group_bin_4380 (RW)
0xda: frame_vm_group_bin_3085 (RW)
0xdb: frame_vm_group_bin_19153 (RW)
0xdc: frame_vm_group_bin_11990 (RW)
0xdd: frame_vm_group_bin_4885 (RW)
0xde: frame_vm_group_bin_20978 (RW)
0xdf: frame_vm_group_bin_13810 (RW)
0xe0: frame_vm_group_bin_6621 (RW)
0xe1: frame_vm_group_bin_22817 (RW)
0xe2: frame_vm_group_bin_15634 (RW)
0xe3: frame_vm_group_bin_8444 (RW)
0xe4: frame_vm_group_bin_1254 (RW)
0xe5: frame_vm_group_bin_21165 (RW)
0xe6: frame_vm_group_bin_10277 (RW)
0xe7: frame_vm_group_bin_3117 (RW)
0xe8: frame_vm_group_bin_19186 (RW)
0xe9: frame_vm_group_bin_15441 (RW)
0xe: frame_vm_group_bin_20476 (RW)
0xea: frame_vm_group_bin_4918 (RW)
0xeb: frame_vm_group_bin_21011 (RW)
0xec: frame_vm_group_bin_13839 (RW)
0xed: frame_vm_group_bin_6654 (RW)
0xee: frame_vm_group_bin_22850 (RW)
0xef: frame_vm_group_bin_15667 (RW)
0xf0: frame_vm_group_bin_8477 (RW)
0xf1: frame_vm_group_bin_1285 (RW)
0xf2: frame_vm_group_bin_2538 (RW)
0xf3: frame_vm_group_bin_10310 (RW)
0xf4: frame_vm_group_bin_3150 (RW)
0xf5: frame_vm_group_bin_19219 (RW)
0xf6: frame_vm_group_bin_20083 (RW)
0xf7: frame_vm_group_bin_4949 (RW)
0xf8: frame_vm_group_bin_21044 (RW)
0xf9: frame_vm_group_bin_13868 (RW)
0xf: frame_vm_group_bin_13279 (RW)
0xfa: frame_vm_group_bin_6688 (RW)
0xfb: frame_vm_group_bin_22884 (RW)
0xfc: frame_vm_group_bin_15701 (RW)
0xfd: frame_vm_group_bin_8511 (RW)
0xfe: frame_vm_group_bin_1318 (RW)
0xff: frame_vm_group_bin_7146 (RW)
}
pt_vm_group_bin_0134 {
0x0: frame_vm_group_bin_9396 (RW)
0x100: frame_vm_group_bin_15421 (RW)
0x101: frame_vm_group_bin_8230 (RW)
0x102: frame_vm_group_bin_2918 (RW)
0x103: frame_vm_group_bin_17266 (RW)
0x104: frame_vm_group_bin_10060 (RW)
0x105: frame_vm_group_bin_2903 (RW)
0x106: frame_vm_group_bin_18973 (RW)
0x107: frame_vm_group_bin_11832 (RW)
0x108: frame_vm_group_bin_4705 (RW)
0x109: frame_vm_group_bin_20827 (RW)
0x10: frame_vm_group_bin_11284 (RW)
0x10a: frame_vm_group_bin_13629 (RW)
0x10b: frame_vm_group_bin_6439 (RW)
0x10c: frame_vm_group_bin_22636 (RW)
0x10d: frame_vm_group_bin_15454 (RW)
0x10e: frame_vm_group_bin_8263 (RW)
0x10f: frame_vm_group_bin_7527 (RW)
0x110: frame_vm_group_bin_17299 (RW)
0x111: frame_vm_group_bin_10093 (RW)
0x112: frame_vm_group_bin_2936 (RW)
0x113: frame_vm_group_bin_19006 (RW)
0x114: frame_vm_group_bin_11860 (RW)
0x115: frame_vm_group_bin_4737 (RW)
0x116: frame_vm_group_bin_20856 (RW)
0x117: frame_vm_group_bin_13661 (RW)
0x118: frame_vm_group_bin_6472 (RW)
0x119: frame_vm_group_bin_22669 (RW)
0x11: frame_vm_group_bin_4099 (RW)
0x11a: frame_vm_group_bin_15488 (RW)
0x11b: frame_vm_group_bin_8296 (RW)
0x11c: frame_vm_group_bin_1108 (RW)
0x11d: frame_vm_group_bin_17333 (RW)
0x11e: frame_vm_group_bin_10127 (RW)
0x11f: frame_vm_group_bin_2970 (RW)
0x120: frame_vm_group_bin_19040 (RW)
0x121: frame_vm_group_bin_5093 (RW)
0x122: frame_vm_group_bin_4771 (RW)
0x123: frame_vm_group_bin_2190 (RW)
0x124: frame_vm_group_bin_13695 (RW)
0x125: frame_vm_group_bin_6506 (RW)
0x126: frame_vm_group_bin_22703 (RW)
0x127: frame_vm_group_bin_15520 (RW)
0x128: frame_vm_group_bin_8329 (RW)
0x129: frame_vm_group_bin_1140 (RW)
0x12: frame_vm_group_bin_20193 (RW)
0x12a: frame_vm_group_bin_17365 (RW)
0x12b: frame_vm_group_bin_10162 (RW)
0x12c: frame_vm_group_bin_3003 (RW)
0x12d: frame_vm_group_bin_19073 (RW)
0x12e: frame_vm_group_bin_11912 (RW)
0x12f: frame_vm_group_bin_4804 (RW)
0x130: frame_vm_group_bin_6824 (RW)
0x131: frame_vm_group_bin_13727 (RW)
0x132: frame_vm_group_bin_6539 (RW)
0x133: frame_vm_group_bin_22736 (RW)
0x134: frame_vm_group_bin_15552 (RW)
0x135: frame_vm_group_bin_8362 (RW)
0x136: frame_vm_group_bin_1173 (RW)
0x137: frame_vm_group_bin_17395 (RW)
0x138: frame_vm_group_bin_10195 (RW)
0x139: frame_vm_group_bin_3036 (RW)
0x13: frame_vm_group_bin_12995 (RW)
0x13a: frame_vm_group_bin_19107 (RW)
0x13b: frame_vm_group_bin_11942 (RW)
0x13c: frame_vm_group_bin_4837 (RW)
0x13d: frame_vm_group_bin_20938 (RW)
0x13e: frame_vm_group_bin_13762 (RW)
0x13f: frame_vm_group_bin_6573 (RW)
0x140: frame_vm_group_bin_22769 (RW)
0x141: frame_vm_group_bin_15586 (RW)
0x142: frame_vm_group_bin_8396 (RW)
0x143: frame_vm_group_bin_1207 (RW)
0x144: frame_vm_group_bin_1458 (RW)
0x145: frame_vm_group_bin_10229 (RW)
0x146: frame_vm_group_bin_3070 (RW)
0x147: frame_vm_group_bin_19138 (RW)
0x148: frame_vm_group_bin_11975 (RW)
0x149: frame_vm_group_bin_4870 (RW)
0x14: frame_vm_group_bin_5877 (RW)
0x14a: frame_vm_group_bin_16215 (RW)
0x14b: frame_vm_group_bin_13795 (RW)
0x14c: frame_vm_group_bin_6606 (RW)
0x14d: frame_vm_group_bin_22802 (RW)
0x14e: frame_vm_group_bin_15619 (RW)
0x14f: frame_vm_group_bin_8429 (RW)
0x150: frame_vm_group_bin_1240 (RW)
0x151: frame_vm_group_bin_6111 (RW)
0x152: frame_vm_group_bin_10262 (RW)
0x153: frame_vm_group_bin_3103 (RW)
0x154: frame_vm_group_bin_19171 (RW)
0x155: frame_vm_group_bin_12007 (RW)
0x156: frame_vm_group_bin_4903 (RW)
0x157: frame_vm_group_bin_20996 (RW)
0x158: frame_vm_group_bin_13826 (RW)
0x159: frame_vm_group_bin_6639 (RW)
0x15: frame_vm_group_bin_22028 (RW)
0x15a: frame_vm_group_bin_22836 (RW)
0x15b: frame_vm_group_bin_15653 (RW)
0x15c: frame_vm_group_bin_8463 (RW)
0x15d: frame_vm_group_bin_12208 (RW)
0x15e: frame_vm_group_bin_17467 (RW)
0x15f: frame_vm_group_bin_10296 (RW)
0x160: frame_vm_group_bin_3136 (RW)
0x161: frame_vm_group_bin_19205 (RW)
0x162: frame_vm_group_bin_12038 (RW)
0x163: frame_vm_group_bin_4935 (RW)
0x164: frame_vm_group_bin_21030 (RW)
0x165: frame_vm_group_bin_0763 (RW)
0x166: frame_vm_group_bin_6673 (RW)
0x167: frame_vm_group_bin_22869 (RW)
0x168: frame_vm_group_bin_15686 (RW)
0x169: frame_vm_group_bin_8496 (RW)
0x16: frame_vm_group_bin_14856 (RW)
0x16a: frame_vm_group_bin_1304 (RW)
0x16b: frame_vm_group_bin_17489 (RW)
0x16c: frame_vm_group_bin_10329 (RW)
0x16d: frame_vm_group_bin_3169 (RW)
0x16e: frame_vm_group_bin_19238 (RW)
0x16f: frame_vm_group_bin_12065 (RW)
0x170: frame_vm_group_bin_4966 (RW)
0x171: frame_vm_group_bin_21064 (RW)
0x172: frame_vm_group_bin_13886 (RW)
0x173: frame_vm_group_bin_6706 (RW)
0x174: frame_vm_group_bin_22902 (RW)
0x175: frame_vm_group_bin_15719 (RW)
0x176: frame_vm_group_bin_8528 (RW)
0x177: frame_vm_group_bin_1336 (RW)
0x178: frame_vm_group_bin_17514 (RW)
0x179: frame_vm_group_bin_10362 (RW)
0x17: frame_vm_group_bin_7641 (RW)
0x17a: frame_vm_group_bin_3203 (RW)
0x17b: frame_vm_group_bin_19272 (RW)
0x17c: frame_vm_group_bin_12099 (RW)
0x17d: frame_vm_group_bin_5000 (RW)
0x17e: frame_vm_group_bin_21098 (RW)
0x17f: frame_vm_group_bin_13920 (RW)
0x180: frame_vm_group_bin_6739 (RW)
0x181: frame_vm_group_bin_22936 (RW)
0x182: frame_vm_group_bin_15753 (RW)
0x183: frame_vm_group_bin_8560 (RW)
0x184: frame_vm_group_bin_1371 (RW)
0x185: frame_vm_group_bin_17541 (RW)
0x186: frame_vm_group_bin_0101 (RW)
0x187: frame_vm_group_bin_3235 (RW)
0x188: frame_vm_group_bin_19305 (RW)
0x189: frame_vm_group_bin_12131 (RW)
0x18: frame_vm_group_bin_0481 (RW)
0x18a: frame_vm_group_bin_5033 (RW)
0x18b: frame_vm_group_bin_21131 (RW)
0x18c: frame_vm_group_bin_13953 (RW)
0x18d: frame_vm_group_bin_6771 (RW)
0x18e: frame_vm_group_bin_22968 (RW)
0x18f: frame_vm_group_bin_15786 (RW)
0x190: frame_vm_group_bin_8593 (RW)
0x191: frame_vm_group_bin_1404 (RW)
0x192: frame_vm_group_bin_17562 (RW)
0x193: frame_vm_group_bin_4765 (RW)
0x194: frame_vm_group_bin_3268 (RW)
0x195: frame_vm_group_bin_19338 (RW)
0x196: frame_vm_group_bin_12163 (RW)
0x197: frame_vm_group_bin_5066 (RW)
0x198: frame_vm_group_bin_21163 (RW)
0x199: frame_vm_group_bin_13986 (RW)
0x19: frame_vm_group_bin_16671 (RW)
0x19a: frame_vm_group_bin_6805 (RW)
0x19b: frame_vm_group_bin_23001 (RW)
0x19c: frame_vm_group_bin_15819 (RW)
0x19d: frame_vm_group_bin_8626 (RW)
0x19e: frame_vm_group_bin_1438 (RW)
0x19f: frame_vm_group_bin_17587 (RW)
0x1: frame_vm_group_bin_2237 (RW)
0x1a0: frame_vm_group_bin_10449 (RW)
0x1a1: frame_vm_group_bin_3302 (RW)
0x1a2: frame_vm_group_bin_19372 (RW)
0x1a3: frame_vm_group_bin_12194 (RW)
0x1a4: frame_vm_group_bin_5101 (RW)
0x1a5: frame_vm_group_bin_21197 (RW)
0x1a6: frame_vm_group_bin_14020 (RW)
0x1a7: frame_vm_group_bin_6835 (RW)
0x1a8: frame_vm_group_bin_23034 (RW)
0x1a9: frame_vm_group_bin_15851 (RW)
0x1a: frame_vm_group_bin_9463 (RW)
0x1aa: frame_vm_group_bin_8659 (RW)
0x1ab: frame_vm_group_bin_1471 (RW)
0x1ac: frame_vm_group_bin_17611 (RW)
0x1ad: frame_vm_group_bin_10482 (RW)
0x1ae: frame_vm_group_bin_3335 (RW)
0x1af: frame_vm_group_bin_19405 (RW)
0x1b0: frame_vm_group_bin_12224 (RW)
0x1b1: frame_vm_group_bin_5134 (RW)
0x1b2: frame_vm_group_bin_21230 (RW)
0x1b3: frame_vm_group_bin_14053 (RW)
0x1b4: frame_vm_group_bin_4058 (RW)
0x1b5: frame_vm_group_bin_23067 (RW)
0x1b6: frame_vm_group_bin_15884 (RW)
0x1b7: frame_vm_group_bin_8693 (RW)
0x1b8: frame_vm_group_bin_1504 (RW)
0x1b9: frame_vm_group_bin_17644 (RW)
0x1b: frame_vm_group_bin_2303 (RW)
0x1ba: frame_vm_group_bin_10516 (RW)
0x1bb: frame_vm_group_bin_3369 (RW)
0x1bc: frame_vm_group_bin_15888 (RW)
0x1bd: frame_vm_group_bin_12257 (RW)
0x1be: frame_vm_group_bin_5168 (RW)
0x1bf: frame_vm_group_bin_21264 (RW)
0x1c0: frame_vm_group_bin_14087 (RW)
0x1c1: frame_vm_group_bin_8696 (RW)
0x1c2: frame_vm_group_bin_23101 (RW)
0x1c3: frame_vm_group_bin_15918 (RW)
0x1c4: frame_vm_group_bin_8727 (RW)
0x1c5: frame_vm_group_bin_1538 (RW)
0x1c6: frame_vm_group_bin_17678 (RW)
0x1c7: frame_vm_group_bin_10548 (RW)
0x1c8: frame_vm_group_bin_3399 (RW)
0x1c9: frame_vm_group_bin_19468 (RW)
0x1c: frame_vm_group_bin_18405 (RW)
0x1ca: frame_vm_group_bin_12290 (RW)
0x1cb: frame_vm_group_bin_5201 (RW)
0x1cc: frame_vm_group_bin_21297 (RW)
0x1cd: frame_vm_group_bin_14120 (RW)
0x1ce: frame_vm_group_bin_6910 (RW)
0x1cf: frame_vm_group_bin_23134 (RW)
0x1d0: frame_vm_group_bin_15951 (RW)
0x1d1: frame_vm_group_bin_8760 (RW)
0x1d2: frame_vm_group_bin_1571 (RW)
0x1d3: frame_vm_group_bin_17704 (RW)
0x1d4: frame_vm_group_bin_10581 (RW)
0x1d5: frame_vm_group_bin_3367 (RW)
0x1d6: frame_vm_group_bin_19501 (RW)
0x1d7: frame_vm_group_bin_12323 (RW)
0x1d8: frame_vm_group_bin_5234 (RW)
0x1d9: frame_vm_group_bin_21328 (RW)
0x1d: frame_vm_group_bin_11318 (RW)
0x1da: frame_vm_group_bin_14154 (RW)
0x1db: frame_vm_group_bin_6942 (RW)
0x1dc: frame_vm_group_bin_23167 (RW)
0x1dd: frame_vm_group_bin_15987 (RW)
0x1de: frame_vm_group_bin_8794 (RW)
0x1df: frame_vm_group_bin_1605 (RW)
0x1e0: frame_vm_group_bin_17732 (RW)
0x1e1: frame_vm_group_bin_10615 (RW)
0x1e2: frame_vm_group_bin_7975 (RW)
0x1e3: frame_vm_group_bin_19535 (RW)
0x1e4: frame_vm_group_bin_12356 (RW)
0x1e5: frame_vm_group_bin_5268 (RW)
0x1e6: frame_vm_group_bin_21362 (RW)
0x1e7: frame_vm_group_bin_14186 (RW)
0x1e8: frame_vm_group_bin_6973 (RW)
0x1e9: frame_vm_group_bin_23199 (RW)
0x1e: frame_vm_group_bin_4132 (RW)
0x1ea: frame_vm_group_bin_16020 (RW)
0x1eb: frame_vm_group_bin_8827 (RW)
0x1ec: frame_vm_group_bin_1638 (RW)
0x1ed: frame_vm_group_bin_17759 (RW)
0x1ee: frame_vm_group_bin_10647 (RW)
0x1ef: frame_vm_group_bin_12631 (RW)
0x1f0: frame_vm_group_bin_19568 (RW)
0x1f1: frame_vm_group_bin_12389 (RW)
0x1f2: frame_vm_group_bin_5301 (RW)
0x1f3: frame_vm_group_bin_21395 (RW)
0x1f4: frame_vm_group_bin_14219 (RW)
0x1f5: frame_vm_group_bin_7006 (RW)
0x1f6: frame_vm_group_bin_23222 (RW)
0x1f7: frame_vm_group_bin_16053 (RW)
0x1f8: frame_vm_group_bin_8860 (RW)
0x1f9: frame_vm_group_bin_1671 (RW)
0x1f: frame_vm_group_bin_20227 (RW)
0x1fa: frame_vm_group_bin_20176 (RW)
0x1fb: frame_vm_group_bin_10680 (RW)
0x1fc: frame_vm_group_bin_3498 (RW)
0x1fd: frame_vm_group_bin_19603 (RW)
0x1fe: frame_vm_group_bin_12423 (RW)
0x1ff: frame_vm_group_bin_5333 (RW)
0x20: frame_vm_group_bin_13031 (RW)
0x21: frame_vm_group_bin_5904 (RW)
0x22: frame_vm_group_bin_21093 (RW)
0x23: frame_vm_group_bin_14890 (RW)
0x24: frame_vm_group_bin_7675 (RW)
0x25: frame_vm_group_bin_0514 (RW)
0x26: frame_vm_group_bin_16704 (RW)
0x27: frame_vm_group_bin_9496 (RW)
0x28: frame_vm_group_bin_2336 (RW)
0x29: frame_vm_group_bin_18437 (RW)
0x2: frame_vm_group_bin_18339 (RW)
0x2a: frame_vm_group_bin_11349 (RW)
0x2b: frame_vm_group_bin_4164 (RW)
0x2c: frame_vm_group_bin_20260 (RW)
0x2d: frame_vm_group_bin_13064 (RW)
0x2e: frame_vm_group_bin_5929 (RW)
0x2f: frame_vm_group_bin_2466 (RW)
0x30: frame_vm_group_bin_14923 (RW)
0x31: frame_vm_group_bin_7708 (RW)
0x32: frame_vm_group_bin_0546 (RW)
0x33: frame_vm_group_bin_16738 (RW)
0x34: frame_vm_group_bin_9529 (RW)
0x35: frame_vm_group_bin_2369 (RW)
0x36: frame_vm_group_bin_18468 (RW)
0x37: frame_vm_group_bin_11381 (RW)
0x38: frame_vm_group_bin_12812 (RW)
0x39: frame_vm_group_bin_20292 (RW)
0x3: frame_vm_group_bin_11251 (RW)
0x3a: frame_vm_group_bin_13098 (RW)
0x3b: frame_vm_group_bin_5951 (RW)
0x3c: frame_vm_group_bin_22106 (RW)
0x3d: frame_vm_group_bin_14957 (RW)
0x3e: frame_vm_group_bin_7741 (RW)
0x3f: frame_vm_group_bin_0578 (RW)
0x40: frame_vm_group_bin_16772 (RW)
0x41: frame_vm_group_bin_9563 (RW)
0x42: frame_vm_group_bin_2403 (RW)
0x43: frame_vm_group_bin_18496 (RW)
0x44: frame_vm_group_bin_11414 (RW)
0x45: frame_vm_group_bin_4230 (RW)
0x46: frame_vm_group_bin_20328 (RW)
0x47: frame_vm_group_bin_13131 (RW)
0x48: frame_vm_group_bin_5978 (RW)
0x49: frame_vm_group_bin_22139 (RW)
0x4: frame_vm_group_bin_4066 (RW)
0x4a: frame_vm_group_bin_14990 (RW)
0x4b: frame_vm_group_bin_7774 (RW)
0x4c: frame_vm_group_bin_0610 (RW)
0x4d: frame_vm_group_bin_16805 (RW)
0x4e: frame_vm_group_bin_9596 (RW)
0x4f: frame_vm_group_bin_2435 (RW)
0x50: frame_vm_group_bin_1740 (RW)
0x51: frame_vm_group_bin_11447 (RW)
0x52: frame_vm_group_bin_4263 (RW)
0x53: frame_vm_group_bin_20361 (RW)
0x54: frame_vm_group_bin_13164 (RW)
0x55: frame_vm_group_bin_6009 (RW)
0x56: frame_vm_group_bin_22172 (RW)
0x57: frame_vm_group_bin_15023 (RW)
0x58: frame_vm_group_bin_7807 (RW)
0x59: frame_vm_group_bin_0642 (RW)
0x5: frame_vm_group_bin_20161 (RW)
0x5a: frame_vm_group_bin_16839 (RW)
0x5b: frame_vm_group_bin_9630 (RW)
0x5c: frame_vm_group_bin_2468 (RW)
0x5d: frame_vm_group_bin_18549 (RW)
0x5e: frame_vm_group_bin_11481 (RW)
0x5f: frame_vm_group_bin_4297 (RW)
0x60: frame_vm_group_bin_20395 (RW)
0x61: frame_vm_group_bin_13198 (RW)
0x62: frame_vm_group_bin_6040 (RW)
0x63: frame_vm_group_bin_22206 (RW)
0x64: frame_vm_group_bin_19664 (RW)
0x65: frame_vm_group_bin_7840 (RW)
0x66: frame_vm_group_bin_0676 (RW)
0x67: frame_vm_group_bin_16871 (RW)
0x68: frame_vm_group_bin_9663 (RW)
0x69: frame_vm_group_bin_2501 (RW)
0x6: frame_vm_group_bin_12962 (RW)
0x6a: frame_vm_group_bin_18578 (RW)
0x6b: frame_vm_group_bin_11514 (RW)
0x6c: frame_vm_group_bin_4330 (RW)
0x6d: frame_vm_group_bin_20428 (RW)
0x6e: frame_vm_group_bin_13231 (RW)
0x6f: frame_vm_group_bin_6063 (RW)
0x70: frame_vm_group_bin_22239 (RW)
0x71: frame_vm_group_bin_1036 (RW)
0x72: frame_vm_group_bin_7873 (RW)
0x73: frame_vm_group_bin_0709 (RW)
0x74: frame_vm_group_bin_16903 (RW)
0x75: frame_vm_group_bin_9695 (RW)
0x76: frame_vm_group_bin_2534 (RW)
0x77: frame_vm_group_bin_18611 (RW)
0x78: frame_vm_group_bin_11547 (RW)
0x79: frame_vm_group_bin_4365 (RW)
0x7: frame_vm_group_bin_5851 (RW)
0x7a: frame_vm_group_bin_20462 (RW)
0x7b: frame_vm_group_bin_13265 (RW)
0x7c: frame_vm_group_bin_6092 (RW)
0x7d: frame_vm_group_bin_22272 (RW)
0x7e: frame_vm_group_bin_15101 (RW)
0x7f: frame_vm_group_bin_7907 (RW)
0x80: frame_vm_group_bin_0743 (RW)
0x81: frame_vm_group_bin_16937 (RW)
0x82: frame_vm_group_bin_9729 (RW)
0x83: frame_vm_group_bin_2568 (RW)
0x84: frame_vm_group_bin_18644 (RW)
0x85: frame_vm_group_bin_18942 (RW)
0x86: frame_vm_group_bin_4399 (RW)
0x87: frame_vm_group_bin_20495 (RW)
0x88: frame_vm_group_bin_13298 (RW)
0x89: frame_vm_group_bin_6123 (RW)
0x8: frame_vm_group_bin_21999 (RW)
0x8a: frame_vm_group_bin_22305 (RW)
0x8b: frame_vm_group_bin_10404 (RW)
0x8c: frame_vm_group_bin_7941 (RW)
0x8d: frame_vm_group_bin_0776 (RW)
0x8e: frame_vm_group_bin_16970 (RW)
0x8f: frame_vm_group_bin_9762 (RW)
0x90: frame_vm_group_bin_2601 (RW)
0x91: frame_vm_group_bin_18677 (RW)
0x92: frame_vm_group_bin_0327 (RW)
0x93: frame_vm_group_bin_4432 (RW)
0x94: frame_vm_group_bin_20528 (RW)
0x95: frame_vm_group_bin_13330 (RW)
0x96: frame_vm_group_bin_6155 (RW)
0x97: frame_vm_group_bin_22338 (RW)
0x98: frame_vm_group_bin_15153 (RW)
0x99: frame_vm_group_bin_7974 (RW)
0x9: frame_vm_group_bin_14823 (RW)
0x9a: frame_vm_group_bin_0809 (RW)
0x9b: frame_vm_group_bin_17004 (RW)
0x9c: frame_vm_group_bin_9796 (RW)
0x9d: frame_vm_group_bin_2635 (RW)
0x9e: frame_vm_group_bin_18710 (RW)
0x9f: frame_vm_group_bin_11628 (RW)
0xa0: frame_vm_group_bin_4466 (RW)
0xa1: frame_vm_group_bin_20562 (RW)
0xa2: frame_vm_group_bin_13364 (RW)
0xa3: frame_vm_group_bin_6188 (RW)
0xa4: frame_vm_group_bin_22371 (RW)
0xa5: frame_vm_group_bin_15187 (RW)
0xa6: frame_vm_group_bin_8006 (RW)
0xa7: frame_vm_group_bin_0842 (RW)
0xa8: frame_vm_group_bin_17037 (RW)
0xa9: frame_vm_group_bin_9829 (RW)
0xa: frame_vm_group_bin_7608 (RW)
0xaa: frame_vm_group_bin_2668 (RW)
0xab: frame_vm_group_bin_18741 (RW)
0xac: frame_vm_group_bin_11650 (RW)
0xad: frame_vm_group_bin_4499 (RW)
0xae: frame_vm_group_bin_20595 (RW)
0xaf: frame_vm_group_bin_13395 (RW)
0xb0: frame_vm_group_bin_6215 (RW)
0xb1: frame_vm_group_bin_22404 (RW)
0xb2: frame_vm_group_bin_15220 (RW)
0xb3: frame_vm_group_bin_8033 (RW)
0xb4: frame_vm_group_bin_0875 (RW)
0xb5: frame_vm_group_bin_17070 (RW)
0xb6: frame_vm_group_bin_9862 (RW)
0xb7: frame_vm_group_bin_2701 (RW)
0xb8: frame_vm_group_bin_18774 (RW)
0xb9: frame_vm_group_bin_11670 (RW)
0xb: frame_vm_group_bin_0448 (RW)
0xba: frame_vm_group_bin_4533 (RW)
0xbb: frame_vm_group_bin_20629 (RW)
0xbc: frame_vm_group_bin_13429 (RW)
0xbd: frame_vm_group_bin_6245 (RW)
0xbe: frame_vm_group_bin_22437 (RW)
0xbf: frame_vm_group_bin_15255 (RW)
0xc0: frame_vm_group_bin_8065 (RW)
0xc1: frame_vm_group_bin_0909 (RW)
0xc2: frame_vm_group_bin_17104 (RW)
0xc3: frame_vm_group_bin_9895 (RW)
0xc4: frame_vm_group_bin_2735 (RW)
0xc5: frame_vm_group_bin_18808 (RW)
0xc6: frame_vm_group_bin_11698 (RW)
0xc7: frame_vm_group_bin_4565 (RW)
0xc8: frame_vm_group_bin_20661 (RW)
0xc9: frame_vm_group_bin_13462 (RW)
0xc: frame_vm_group_bin_16638 (RW)
0xca: frame_vm_group_bin_6277 (RW)
0xcb: frame_vm_group_bin_22470 (RW)
0xcc: frame_vm_group_bin_15287 (RW)
0xcd: frame_vm_group_bin_8097 (RW)
0xce: frame_vm_group_bin_0942 (RW)
0xcf: frame_vm_group_bin_17137 (RW)
0xd0: frame_vm_group_bin_9928 (RW)
0xd1: frame_vm_group_bin_2768 (RW)
0xd2: frame_vm_group_bin_18842 (RW)
0xd3: frame_vm_group_bin_11725 (RW)
0xd4: frame_vm_group_bin_22246 (RW)
0xd5: frame_vm_group_bin_20694 (RW)
0xd6: frame_vm_group_bin_13495 (RW)
0xd7: frame_vm_group_bin_6310 (RW)
0xd8: frame_vm_group_bin_22503 (RW)
0xd9: frame_vm_group_bin_15320 (RW)
0xd: frame_vm_group_bin_9429 (RW)
0xda: frame_vm_group_bin_8130 (RW)
0xdb: frame_vm_group_bin_0976 (RW)
0xdc: frame_vm_group_bin_10795 (RW)
0xdd: frame_vm_group_bin_9960 (RW)
0xde: frame_vm_group_bin_2802 (RW)
0xdf: frame_vm_group_bin_18876 (RW)
0xe0: frame_vm_group_bin_11748 (RW)
0xe1: frame_vm_group_bin_3609 (RW)
0xe2: frame_vm_group_bin_20728 (RW)
0xe3: frame_vm_group_bin_13529 (RW)
0xe4: frame_vm_group_bin_6343 (RW)
0xe5: frame_vm_group_bin_22536 (RW)
0xe6: frame_vm_group_bin_15354 (RW)
0xe7: frame_vm_group_bin_8163 (RW)
0xe8: frame_vm_group_bin_1009 (RW)
0xe9: frame_vm_group_bin_17200 (RW)
0xe: frame_vm_group_bin_2269 (RW)
0xea: frame_vm_group_bin_9993 (RW)
0xeb: frame_vm_group_bin_2835 (RW)
0xec: frame_vm_group_bin_18909 (RW)
0xed: frame_vm_group_bin_11771 (RW)
0xee: frame_vm_group_bin_4640 (RW)
0xef: frame_vm_group_bin_20761 (RW)
0xf0: frame_vm_group_bin_13562 (RW)
0xf1: frame_vm_group_bin_6375 (RW)
0xf2: frame_vm_group_bin_22569 (RW)
0xf3: frame_vm_group_bin_15387 (RW)
0xf4: frame_vm_group_bin_8196 (RW)
0xf5: frame_vm_group_bin_21538 (RW)
0xf6: frame_vm_group_bin_17233 (RW)
0xf7: frame_vm_group_bin_10026 (RW)
0xf8: frame_vm_group_bin_2867 (RW)
0xf9: frame_vm_group_bin_15816 (RW)
0xf: frame_vm_group_bin_18372 (RW)
0xfa: frame_vm_group_bin_11799 (RW)
0xfb: frame_vm_group_bin_4674 (RW)
0xfc: frame_vm_group_bin_20795 (RW)
0xfd: frame_vm_group_bin_13596 (RW)
0xfe: frame_vm_group_bin_6406 (RW)
0xff: frame_vm_group_bin_22603 (RW)
}
pt_vm_group_bin_0167 {
0x0: frame_vm_group_bin_19948 (RW)
0x100: frame_vm_group_bin_2685 (RW)
0x101: frame_vm_group_bin_18758 (RW)
0x102: frame_vm_group_bin_11660 (RW)
0x103: frame_vm_group_bin_4516 (RW)
0x104: frame_vm_group_bin_20612 (RW)
0x105: frame_vm_group_bin_13412 (RW)
0x106: frame_vm_group_bin_6230 (RW)
0x107: frame_vm_group_bin_22420 (RW)
0x108: frame_vm_group_bin_15238 (RW)
0x109: frame_vm_group_bin_8049 (RW)
0x10: frame_vm_group_bin_21816 (RW)
0x10a: frame_vm_group_bin_0892 (RW)
0x10b: frame_vm_group_bin_17087 (RW)
0x10c: frame_vm_group_bin_9879 (RW)
0x10d: frame_vm_group_bin_2718 (RW)
0x10e: frame_vm_group_bin_18791 (RW)
0x10f: frame_vm_group_bin_11684 (RW)
0x110: frame_vm_group_bin_4549 (RW)
0x111: frame_vm_group_bin_20645 (RW)
0x112: frame_vm_group_bin_13445 (RW)
0x113: frame_vm_group_bin_6261 (RW)
0x114: frame_vm_group_bin_22453 (RW)
0x115: frame_vm_group_bin_15271 (RW)
0x116: frame_vm_group_bin_8081 (RW)
0x117: frame_vm_group_bin_0925 (RW)
0x118: frame_vm_group_bin_17120 (RW)
0x119: frame_vm_group_bin_9911 (RW)
0x11: frame_vm_group_bin_14641 (RW)
0x11a: frame_vm_group_bin_2752 (RW)
0x11b: frame_vm_group_bin_18827 (RW)
0x11c: frame_vm_group_bin_11713 (RW)
0x11d: frame_vm_group_bin_4578 (RW)
0x11e: frame_vm_group_bin_20678 (RW)
0x11f: frame_vm_group_bin_13479 (RW)
0x120: frame_vm_group_bin_6294 (RW)
0x121: frame_vm_group_bin_22487 (RW)
0x122: frame_vm_group_bin_15304 (RW)
0x123: frame_vm_group_bin_8113 (RW)
0x124: frame_vm_group_bin_0959 (RW)
0x125: frame_vm_group_bin_17153 (RW)
0x126: frame_vm_group_bin_9943 (RW)
0x127: frame_vm_group_bin_2785 (RW)
0x128: frame_vm_group_bin_18859 (RW)
0x129: frame_vm_group_bin_11737 (RW)
0x12: frame_vm_group_bin_7427 (RW)
0x12a: frame_vm_group_bin_3820 (RW)
0x12b: frame_vm_group_bin_20711 (RW)
0x12c: frame_vm_group_bin_13512 (RW)
0x12d: frame_vm_group_bin_6326 (RW)
0x12e: frame_vm_group_bin_22520 (RW)
0x12f: frame_vm_group_bin_15337 (RW)
0x130: frame_vm_group_bin_8146 (RW)
0x131: frame_vm_group_bin_0992 (RW)
0x132: frame_vm_group_bin_17185 (RW)
0x133: frame_vm_group_bin_9976 (RW)
0x134: frame_vm_group_bin_2818 (RW)
0x135: frame_vm_group_bin_18892 (RW)
0x136: frame_vm_group_bin_11758 (RW)
0x137: frame_vm_group_bin_4625 (RW)
0x138: frame_vm_group_bin_20744 (RW)
0x139: frame_vm_group_bin_13545 (RW)
0x13: frame_vm_group_bin_0277 (RW)
0x13a: frame_vm_group_bin_6360 (RW)
0x13b: frame_vm_group_bin_22553 (RW)
0x13c: frame_vm_group_bin_15371 (RW)
0x13d: frame_vm_group_bin_8180 (RW)
0x13e: frame_vm_group_bin_1023 (RW)
0x13f: frame_vm_group_bin_17217 (RW)
0x140: frame_vm_group_bin_10010 (RW)
0x141: frame_vm_group_bin_2852 (RW)
0x142: frame_vm_group_bin_18926 (RW)
0x143: frame_vm_group_bin_11784 (RW)
0x144: frame_vm_group_bin_4657 (RW)
0x145: frame_vm_group_bin_20778 (RW)
0x146: frame_vm_group_bin_13579 (RW)
0x147: frame_vm_group_bin_6390 (RW)
0x148: frame_vm_group_bin_22586 (RW)
0x149: frame_vm_group_bin_15404 (RW)
0x14: frame_vm_group_bin_16456 (RW)
0x14a: frame_vm_group_bin_8213 (RW)
0x14b: frame_vm_group_bin_3131 (RW)
0x14c: frame_vm_group_bin_17249 (RW)
0x14d: frame_vm_group_bin_10043 (RW)
0x14e: frame_vm_group_bin_2886 (RW)
0x14f: frame_vm_group_bin_18958 (RW)
0x150: frame_vm_group_bin_11815 (RW)
0x151: frame_vm_group_bin_4689 (RW)
0x152: frame_vm_group_bin_20811 (RW)
0x153: frame_vm_group_bin_13612 (RW)
0x154: frame_vm_group_bin_6422 (RW)
0x155: frame_vm_group_bin_22619 (RW)
0x156: frame_vm_group_bin_15437 (RW)
0x157: frame_vm_group_bin_8246 (RW)
0x158: frame_vm_group_bin_1066 (RW)
0x159: frame_vm_group_bin_17282 (RW)
0x15: frame_vm_group_bin_4812 (RW)
0x15a: frame_vm_group_bin_10077 (RW)
0x15b: frame_vm_group_bin_2920 (RW)
0x15c: frame_vm_group_bin_18990 (RW)
0x15d: frame_vm_group_bin_11846 (RW)
0x15e: frame_vm_group_bin_4721 (RW)
0x15f: frame_vm_group_bin_20844 (RW)
0x160: frame_vm_group_bin_13645 (RW)
0x161: frame_vm_group_bin_6456 (RW)
0x162: frame_vm_group_bin_22653 (RW)
0x163: frame_vm_group_bin_15471 (RW)
0x164: frame_vm_group_bin_8279 (RW)
0x165: frame_vm_group_bin_12395 (RW)
0x166: frame_vm_group_bin_17316 (RW)
0x167: frame_vm_group_bin_10110 (RW)
0x168: frame_vm_group_bin_2953 (RW)
0x169: frame_vm_group_bin_19023 (RW)
0x16: frame_vm_group_bin_2093 (RW)
0x16a: frame_vm_group_bin_11875 (RW)
0x16b: frame_vm_group_bin_4754 (RW)
0x16c: frame_vm_group_bin_2397 (RW)
0x16d: frame_vm_group_bin_13678 (RW)
0x16e: frame_vm_group_bin_6489 (RW)
0x16f: frame_vm_group_bin_22686 (RW)
0x170: frame_vm_group_bin_15504 (RW)
0x171: frame_vm_group_bin_8312 (RW)
0x172: frame_vm_group_bin_1123 (RW)
0x173: frame_vm_group_bin_17349 (RW)
0x174: frame_vm_group_bin_10143 (RW)
0x175: frame_vm_group_bin_2986 (RW)
0x176: frame_vm_group_bin_19056 (RW)
0x177: frame_vm_group_bin_11898 (RW)
0x178: frame_vm_group_bin_4787 (RW)
0x179: frame_vm_group_bin_20895 (RW)
0x17: frame_vm_group_bin_18189 (RW)
0x17a: frame_vm_group_bin_5677 (RW)
0x17b: frame_vm_group_bin_6523 (RW)
0x17c: frame_vm_group_bin_22720 (RW)
0x17d: frame_vm_group_bin_15537 (RW)
0x17e: frame_vm_group_bin_8346 (RW)
0x17f: frame_vm_group_bin_1157 (RW)
0x180: frame_vm_group_bin_17382 (RW)
0x181: frame_vm_group_bin_10179 (RW)
0x182: frame_vm_group_bin_3020 (RW)
0x183: frame_vm_group_bin_19090 (RW)
0x184: frame_vm_group_bin_11928 (RW)
0x185: frame_vm_group_bin_4820 (RW)
0x186: frame_vm_group_bin_11729 (RW)
0x187: frame_vm_group_bin_13744 (RW)
0x188: frame_vm_group_bin_6556 (RW)
0x189: frame_vm_group_bin_22752 (RW)
0x18: frame_vm_group_bin_11101 (RW)
0x18a: frame_vm_group_bin_15569 (RW)
0x18b: frame_vm_group_bin_8379 (RW)
0x18c: frame_vm_group_bin_1190 (RW)
0x18d: frame_vm_group_bin_10148 (RW)
0x18e: frame_vm_group_bin_10212 (RW)
0x18f: frame_vm_group_bin_3053 (RW)
0x190: frame_vm_group_bin_19122 (RW)
0x191: frame_vm_group_bin_11958 (RW)
0x192: frame_vm_group_bin_4853 (RW)
0x193: frame_vm_group_bin_16412 (RW)
0x194: frame_vm_group_bin_13778 (RW)
0x195: frame_vm_group_bin_6589 (RW)
0x196: frame_vm_group_bin_22785 (RW)
0x197: frame_vm_group_bin_15602 (RW)
0x198: frame_vm_group_bin_8412 (RW)
0x199: frame_vm_group_bin_1223 (RW)
0x19: frame_vm_group_bin_3916 (RW)
0x19a: frame_vm_group_bin_17435 (RW)
0x19b: frame_vm_group_bin_10246 (RW)
0x19c: frame_vm_group_bin_3087 (RW)
0x19d: frame_vm_group_bin_19155 (RW)
0x19e: frame_vm_group_bin_11991 (RW)
0x19f: frame_vm_group_bin_4887 (RW)
0x1: frame_vm_group_bin_12747 (RW)
0x1a0: frame_vm_group_bin_20980 (RW)
0x1a1: frame_vm_group_bin_13812 (RW)
0x1a2: frame_vm_group_bin_6623 (RW)
0x1a3: frame_vm_group_bin_22819 (RW)
0x1a4: frame_vm_group_bin_15636 (RW)
0x1a5: frame_vm_group_bin_8446 (RW)
0x1a6: frame_vm_group_bin_1256 (RW)
0x1a7: frame_vm_group_bin_11055 (RW)
0x1a8: frame_vm_group_bin_10279 (RW)
0x1a9: frame_vm_group_bin_3119 (RW)
0x1a: frame_vm_group_bin_20013 (RW)
0x1aa: frame_vm_group_bin_19188 (RW)
0x1ab: frame_vm_group_bin_12022 (RW)
0x1ac: frame_vm_group_bin_4920 (RW)
0x1ad: frame_vm_group_bin_21013 (RW)
0x1ae: frame_vm_group_bin_13841 (RW)
0x1af: frame_vm_group_bin_6656 (RW)
0x1b0: frame_vm_group_bin_22852 (RW)
0x1b1: frame_vm_group_bin_15669 (RW)
0x1b2: frame_vm_group_bin_8479 (RW)
0x1b3: frame_vm_group_bin_1287 (RW)
0x1b4: frame_vm_group_bin_17477 (RW)
0x1b5: frame_vm_group_bin_10312 (RW)
0x1b6: frame_vm_group_bin_3152 (RW)
0x1b7: frame_vm_group_bin_19221 (RW)
0x1b8: frame_vm_group_bin_12051 (RW)
0x1b9: frame_vm_group_bin_4951 (RW)
0x1b: frame_vm_group_bin_12814 (RW)
0x1ba: frame_vm_group_bin_21048 (RW)
0x1bb: frame_vm_group_bin_13871 (RW)
0x1bc: frame_vm_group_bin_6690 (RW)
0x1bd: frame_vm_group_bin_22886 (RW)
0x1be: frame_vm_group_bin_15703 (RW)
0x1bf: frame_vm_group_bin_8512 (RW)
0x1c0: frame_vm_group_bin_1320 (RW)
0x1c1: frame_vm_group_bin_17500 (RW)
0x1c2: frame_vm_group_bin_10346 (RW)
0x1c3: frame_vm_group_bin_3186 (RW)
0x1c4: frame_vm_group_bin_19255 (RW)
0x1c5: frame_vm_group_bin_12082 (RW)
0x1c6: frame_vm_group_bin_4983 (RW)
0x1c7: frame_vm_group_bin_21081 (RW)
0x1c8: frame_vm_group_bin_13903 (RW)
0x1c9: frame_vm_group_bin_6722 (RW)
0x1c: frame_vm_group_bin_5747 (RW)
0x1ca: frame_vm_group_bin_22919 (RW)
0x1cb: frame_vm_group_bin_15736 (RW)
0x1cc: frame_vm_group_bin_8545 (RW)
0x1cd: frame_vm_group_bin_1353 (RW)
0x1ce: frame_vm_group_bin_17528 (RW)
0x1cf: frame_vm_group_bin_10379 (RW)
0x1d0: frame_vm_group_bin_3219 (RW)
0x1d1: frame_vm_group_bin_19288 (RW)
0x1d2: frame_vm_group_bin_12114 (RW)
0x1d3: frame_vm_group_bin_5016 (RW)
0x1d4: frame_vm_group_bin_21114 (RW)
0x1d5: frame_vm_group_bin_13936 (RW)
0x1d6: frame_vm_group_bin_6755 (RW)
0x1d7: frame_vm_group_bin_22952 (RW)
0x1d8: frame_vm_group_bin_15769 (RW)
0x1d9: frame_vm_group_bin_8576 (RW)
0x1d: frame_vm_group_bin_21850 (RW)
0x1da: frame_vm_group_bin_1388 (RW)
0x1db: frame_vm_group_bin_17553 (RW)
0x1dc: frame_vm_group_bin_10406 (RW)
0x1dd: frame_vm_group_bin_3252 (RW)
0x1de: frame_vm_group_bin_19322 (RW)
0x1df: frame_vm_group_bin_12148 (RW)
0x1e0: frame_vm_group_bin_5050 (RW)
0x1e1: frame_vm_group_bin_21147 (RW)
0x1e2: frame_vm_group_bin_13970 (RW)
0x1e3: frame_vm_group_bin_6788 (RW)
0x1e4: frame_vm_group_bin_22985 (RW)
0x1e5: frame_vm_group_bin_15802 (RW)
0x1e6: frame_vm_group_bin_8609 (RW)
0x1e7: frame_vm_group_bin_1421 (RW)
0x1e8: frame_vm_group_bin_17574 (RW)
0x1e9: frame_vm_group_bin_9605 (RW)
0x1e: frame_vm_group_bin_14675 (RW)
0x1ea: frame_vm_group_bin_3285 (RW)
0x1eb: frame_vm_group_bin_19355 (RW)
0x1ec: frame_vm_group_bin_12178 (RW)
0x1ed: frame_vm_group_bin_5084 (RW)
0x1ee: frame_vm_group_bin_21180 (RW)
0x1ef: frame_vm_group_bin_14003 (RW)
0x1f0: frame_vm_group_bin_6819 (RW)
0x1f1: frame_vm_group_bin_23017 (RW)
0x1f2: frame_vm_group_bin_15834 (RW)
0x1f3: frame_vm_group_bin_8642 (RW)
0x1f4: frame_vm_group_bin_1454 (RW)
0x1f5: frame_vm_group_bin_17597 (RW)
0x1f6: frame_vm_group_bin_10465 (RW)
0x1f7: frame_vm_group_bin_3318 (RW)
0x1f8: frame_vm_group_bin_19388 (RW)
0x1f9: frame_vm_group_bin_12207 (RW)
0x1f: frame_vm_group_bin_7461 (RW)
0x1fa: frame_vm_group_bin_5118 (RW)
0x1fb: frame_vm_group_bin_21214 (RW)
0x1fc: frame_vm_group_bin_14037 (RW)
0x1fd: frame_vm_group_bin_6848 (RW)
0x1fe: frame_vm_group_bin_23051 (RW)
0x1ff: frame_vm_group_bin_15868 (RW)
0x20: frame_vm_group_bin_0308 (RW)
0x21: frame_vm_group_bin_16490 (RW)
0x22: frame_vm_group_bin_9439 (RW)
0x23: frame_vm_group_bin_2128 (RW)
0x24: frame_vm_group_bin_18222 (RW)
0x25: frame_vm_group_bin_11134 (RW)
0x26: frame_vm_group_bin_3949 (RW)
0x27: frame_vm_group_bin_20046 (RW)
0x28: frame_vm_group_bin_12846 (RW)
0x29: frame_vm_group_bin_22740 (RW)
0x2: frame_vm_group_bin_5683 (RW)
0x2a: frame_vm_group_bin_21883 (RW)
0x2b: frame_vm_group_bin_14708 (RW)
0x2c: frame_vm_group_bin_7494 (RW)
0x2d: frame_vm_group_bin_0340 (RW)
0x2e: frame_vm_group_bin_16523 (RW)
0x2f: frame_vm_group_bin_14107 (RW)
0x30: frame_vm_group_bin_2161 (RW)
0x31: frame_vm_group_bin_18255 (RW)
0x32: frame_vm_group_bin_11167 (RW)
0x33: frame_vm_group_bin_3982 (RW)
0x34: frame_vm_group_bin_20079 (RW)
0x35: frame_vm_group_bin_12879 (RW)
0x36: frame_vm_group_bin_4105 (RW)
0x37: frame_vm_group_bin_21916 (RW)
0x38: frame_vm_group_bin_14740 (RW)
0x39: frame_vm_group_bin_7526 (RW)
0x3: frame_vm_group_bin_21782 (RW)
0x3a: frame_vm_group_bin_0372 (RW)
0x3b: frame_vm_group_bin_16556 (RW)
0x3c: frame_vm_group_bin_9345 (RW)
0x3d: frame_vm_group_bin_2194 (RW)
0x3e: frame_vm_group_bin_18289 (RW)
0x3f: frame_vm_group_bin_11201 (RW)
0x40: frame_vm_group_bin_4016 (RW)
0x41: frame_vm_group_bin_20112 (RW)
0x42: frame_vm_group_bin_12913 (RW)
0x43: frame_vm_group_bin_5814 (RW)
0x44: frame_vm_group_bin_21949 (RW)
0x45: frame_vm_group_bin_14774 (RW)
0x46: frame_vm_group_bin_7558 (RW)
0x47: frame_vm_group_bin_0402 (RW)
0x48: frame_vm_group_bin_16589 (RW)
0x49: frame_vm_group_bin_9378 (RW)
0x4: frame_vm_group_bin_14608 (RW)
0x4a: frame_vm_group_bin_22030 (RW)
0x4b: frame_vm_group_bin_18322 (RW)
0x4c: frame_vm_group_bin_11234 (RW)
0x4d: frame_vm_group_bin_4049 (RW)
0x4e: frame_vm_group_bin_20145 (RW)
0x4f: frame_vm_group_bin_12945 (RW)
0x50: frame_vm_group_bin_5839 (RW)
0x51: frame_vm_group_bin_21982 (RW)
0x52: frame_vm_group_bin_14806 (RW)
0x53: frame_vm_group_bin_7591 (RW)
0x54: frame_vm_group_bin_0431 (RW)
0x55: frame_vm_group_bin_16621 (RW)
0x56: frame_vm_group_bin_9412 (RW)
0x57: frame_vm_group_bin_2252 (RW)
0x58: frame_vm_group_bin_18355 (RW)
0x59: frame_vm_group_bin_11267 (RW)
0x5: frame_vm_group_bin_7394 (RW)
0x5a: frame_vm_group_bin_4083 (RW)
0x5b: frame_vm_group_bin_20178 (RW)
0x5c: frame_vm_group_bin_12979 (RW)
0x5d: frame_vm_group_bin_5863 (RW)
0x5e: frame_vm_group_bin_22015 (RW)
0x5f: frame_vm_group_bin_14840 (RW)
0x60: frame_vm_group_bin_7625 (RW)
0x61: frame_vm_group_bin_0465 (RW)
0x62: frame_vm_group_bin_16655 (RW)
0x63: frame_vm_group_bin_9446 (RW)
0x64: frame_vm_group_bin_2286 (RW)
0x65: frame_vm_group_bin_18389 (RW)
0x66: frame_vm_group_bin_11301 (RW)
0x67: frame_vm_group_bin_4115 (RW)
0x68: frame_vm_group_bin_20210 (RW)
0x69: frame_vm_group_bin_13014 (RW)
0x6: frame_vm_group_bin_0253 (RW)
0x6a: frame_vm_group_bin_5889 (RW)
0x6b: frame_vm_group_bin_1362 (RW)
0x6c: frame_vm_group_bin_14873 (RW)
0x6d: frame_vm_group_bin_7658 (RW)
0x6e: frame_vm_group_bin_0497 (RW)
0x6f: frame_vm_group_bin_16688 (RW)
0x70: frame_vm_group_bin_9479 (RW)
0x71: frame_vm_group_bin_2319 (RW)
0x72: frame_vm_group_bin_18420 (RW)
0x73: frame_vm_group_bin_11334 (RW)
0x74: frame_vm_group_bin_4148 (RW)
0x75: frame_vm_group_bin_20243 (RW)
0x76: frame_vm_group_bin_13047 (RW)
0x77: frame_vm_group_bin_5915 (RW)
0x78: frame_vm_group_bin_22061 (RW)
0x79: frame_vm_group_bin_14906 (RW)
0x7: frame_vm_group_bin_16423 (RW)
0x7a: frame_vm_group_bin_7692 (RW)
0x7b: frame_vm_group_bin_0530 (RW)
0x7c: frame_vm_group_bin_16722 (RW)
0x7d: frame_vm_group_bin_9513 (RW)
0x7e: frame_vm_group_bin_2353 (RW)
0x7f: frame_vm_group_bin_18454 (RW)
0x80: frame_vm_group_bin_11366 (RW)
0x81: frame_vm_group_bin_4181 (RW)
0x82: frame_vm_group_bin_20276 (RW)
0x83: frame_vm_group_bin_13081 (RW)
0x84: frame_vm_group_bin_5939 (RW)
0x85: frame_vm_group_bin_22090 (RW)
0x86: frame_vm_group_bin_14940 (RW)
0x87: frame_vm_group_bin_7724 (RW)
0x88: frame_vm_group_bin_0561 (RW)
0x89: frame_vm_group_bin_16755 (RW)
0x8: frame_vm_group_bin_0133 (RW)
0x8a: frame_vm_group_bin_9546 (RW)
0x8b: frame_vm_group_bin_2386 (RW)
0x8c: frame_vm_group_bin_18482 (RW)
0x8d: frame_vm_group_bin_11398 (RW)
0x8e: frame_vm_group_bin_4213 (RW)
0x8f: frame_vm_group_bin_20309 (RW)
0x90: frame_vm_group_bin_13114 (RW)
0x91: frame_vm_group_bin_5964 (RW)
0x92: frame_vm_group_bin_22122 (RW)
0x93: frame_vm_group_bin_14973 (RW)
0x94: frame_vm_group_bin_7757 (RW)
0x95: frame_vm_group_bin_0593 (RW)
0x96: frame_vm_group_bin_16788 (RW)
0x97: frame_vm_group_bin_9579 (RW)
0x98: frame_vm_group_bin_2419 (RW)
0x99: frame_vm_group_bin_18509 (RW)
0x9: frame_vm_group_bin_2060 (RW)
0x9a: frame_vm_group_bin_11431 (RW)
0x9b: frame_vm_group_bin_4247 (RW)
0x9c: frame_vm_group_bin_20345 (RW)
0x9d: frame_vm_group_bin_13148 (RW)
0x9e: frame_vm_group_bin_5993 (RW)
0x9f: frame_vm_group_bin_22156 (RW)
0xa0: frame_vm_group_bin_15007 (RW)
0xa1: frame_vm_group_bin_7791 (RW)
0xa2: frame_vm_group_bin_0625 (RW)
0xa3: frame_vm_group_bin_16822 (RW)
0xa4: frame_vm_group_bin_9613 (RW)
0xa5: frame_vm_group_bin_2452 (RW)
0xa6: frame_vm_group_bin_6593 (RW)
0xa7: frame_vm_group_bin_11464 (RW)
0xa8: frame_vm_group_bin_4280 (RW)
0xa9: frame_vm_group_bin_20378 (RW)
0xa: frame_vm_group_bin_18156 (RW)
0xaa: frame_vm_group_bin_13181 (RW)
0xab: frame_vm_group_bin_6024 (RW)
0xac: frame_vm_group_bin_22189 (RW)
0xad: frame_vm_group_bin_15038 (RW)
0xae: frame_vm_group_bin_7824 (RW)
0xaf: frame_vm_group_bin_0659 (RW)
0xb0: frame_vm_group_bin_16855 (RW)
0xb1: frame_vm_group_bin_9646 (RW)
0xb2: frame_vm_group_bin_2484 (RW)
0xb3: frame_vm_group_bin_11338 (RW)
0xb4: frame_vm_group_bin_11497 (RW)
0xb5: frame_vm_group_bin_4313 (RW)
0xb6: frame_vm_group_bin_20411 (RW)
0xb7: frame_vm_group_bin_13214 (RW)
0xb8: frame_vm_group_bin_6050 (RW)
0xb9: frame_vm_group_bin_22222 (RW)
0xb: frame_vm_group_bin_11068 (RW)
0xba: frame_vm_group_bin_15063 (RW)
0xbb: frame_vm_group_bin_7857 (RW)
0xbc: frame_vm_group_bin_0693 (RW)
0xbd: frame_vm_group_bin_16888 (RW)
0xbe: frame_vm_group_bin_18776 (RW)
0xbf: frame_vm_group_bin_2518 (RW)
0xc0: frame_vm_group_bin_18595 (RW)
0xc1: frame_vm_group_bin_11531 (RW)
0xc2: frame_vm_group_bin_4349 (RW)
0xc3: frame_vm_group_bin_20445 (RW)
0xc4: frame_vm_group_bin_13248 (RW)
0xc5: frame_vm_group_bin_6076 (RW)
0xc6: frame_vm_group_bin_22256 (RW)
0xc7: frame_vm_group_bin_5918 (RW)
0xc8: frame_vm_group_bin_7890 (RW)
0xc9: frame_vm_group_bin_0726 (RW)
0xc: frame_vm_group_bin_3883 (RW)
0xca: frame_vm_group_bin_16920 (RW)
0xcb: frame_vm_group_bin_9712 (RW)
0xcc: frame_vm_group_bin_2551 (RW)
0xcd: frame_vm_group_bin_18628 (RW)
0xce: frame_vm_group_bin_11562 (RW)
0xcf: frame_vm_group_bin_4382 (RW)
0xd0: frame_vm_group_bin_20478 (RW)
0xd1: frame_vm_group_bin_13281 (RW)
0xd2: frame_vm_group_bin_6107 (RW)
0xd3: frame_vm_group_bin_22288 (RW)
0xd4: frame_vm_group_bin_15114 (RW)
0xd5: frame_vm_group_bin_7923 (RW)
0xd6: frame_vm_group_bin_0759 (RW)
0xd7: frame_vm_group_bin_16953 (RW)
0xd8: frame_vm_group_bin_9745 (RW)
0xd9: frame_vm_group_bin_2584 (RW)
0xd: frame_vm_group_bin_19981 (RW)
0xda: frame_vm_group_bin_18661 (RW)
0xdb: frame_vm_group_bin_11590 (RW)
0xdc: frame_vm_group_bin_4416 (RW)
0xdd: frame_vm_group_bin_20512 (RW)
0xde: frame_vm_group_bin_13315 (RW)
0xdf: frame_vm_group_bin_18074 (RW)
0xe0: frame_vm_group_bin_22322 (RW)
0xe1: frame_vm_group_bin_15250 (RW)
0xe2: frame_vm_group_bin_7958 (RW)
0xe3: frame_vm_group_bin_0793 (RW)
0xe4: frame_vm_group_bin_16987 (RW)
0xe5: frame_vm_group_bin_9779 (RW)
0xe6: frame_vm_group_bin_2618 (RW)
0xe7: frame_vm_group_bin_18694 (RW)
0xe8: frame_vm_group_bin_5259 (RW)
0xe9: frame_vm_group_bin_4449 (RW)
0xe: frame_vm_group_bin_12780 (RW)
0xea: frame_vm_group_bin_20545 (RW)
0xeb: frame_vm_group_bin_13347 (RW)
0xec: frame_vm_group_bin_6172 (RW)
0xed: frame_vm_group_bin_22354 (RW)
0xee: frame_vm_group_bin_15170 (RW)
0xef: frame_vm_group_bin_7990 (RW)
0xf0: frame_vm_group_bin_0825 (RW)
0xf1: frame_vm_group_bin_17020 (RW)
0xf2: frame_vm_group_bin_9812 (RW)
0xf3: frame_vm_group_bin_2651 (RW)
0xf4: frame_vm_group_bin_18726 (RW)
0xf5: frame_vm_group_bin_11637 (RW)
0xf6: frame_vm_group_bin_4482 (RW)
0xf7: frame_vm_group_bin_20578 (RW)
0xf8: frame_vm_group_bin_5628 (RW)
0xf9: frame_vm_group_bin_6203 (RW)
0xf: frame_vm_group_bin_5716 (RW)
0xfa: frame_vm_group_bin_22388 (RW)
0xfb: frame_vm_group_bin_15204 (RW)
0xfc: frame_vm_group_bin_8021 (RW)
0xfd: frame_vm_group_bin_0859 (RW)
0xfe: frame_vm_group_bin_17054 (RW)
0xff: frame_vm_group_bin_9846 (RW)
}
pt_vm_group_bin_0176 {
0x0: frame_vm_group_bin_10895 (RW)
0x100: frame_vm_group_bin_16913 (RW)
0x101: frame_vm_group_bin_9705 (RW)
0x102: frame_vm_group_bin_2544 (RW)
0x103: frame_vm_group_bin_18621 (RW)
0x104: frame_vm_group_bin_11557 (RW)
0x105: frame_vm_group_bin_4375 (RW)
0x106: frame_vm_group_bin_20471 (RW)
0x107: frame_vm_group_bin_13274 (RW)
0x108: frame_vm_group_bin_6101 (RW)
0x109: frame_vm_group_bin_22281 (RW)
0x10: frame_vm_group_bin_0281 (RW)
0x10a: frame_vm_group_bin_14742 (RW)
0x10b: frame_vm_group_bin_7916 (RW)
0x10c: frame_vm_group_bin_0752 (RW)
0x10d: frame_vm_group_bin_16946 (RW)
0x10e: frame_vm_group_bin_9738 (RW)
0x10f: frame_vm_group_bin_2577 (RW)
0x110: frame_vm_group_bin_18653 (RW)
0x111: frame_vm_group_bin_4717 (RW)
0x112: frame_vm_group_bin_4408 (RW)
0x113: frame_vm_group_bin_20504 (RW)
0x114: frame_vm_group_bin_13307 (RW)
0x115: frame_vm_group_bin_6132 (RW)
0x116: frame_vm_group_bin_22314 (RW)
0x117: frame_vm_group_bin_19366 (RW)
0x118: frame_vm_group_bin_7950 (RW)
0x119: frame_vm_group_bin_0785 (RW)
0x11: frame_vm_group_bin_5578 (RW)
0x11a: frame_vm_group_bin_16980 (RW)
0x11b: frame_vm_group_bin_9772 (RW)
0x11c: frame_vm_group_bin_2611 (RW)
0x11d: frame_vm_group_bin_18687 (RW)
0x11e: frame_vm_group_bin_11610 (RW)
0x11f: frame_vm_group_bin_4442 (RW)
0x120: frame_vm_group_bin_20538 (RW)
0x121: frame_vm_group_bin_13340 (RW)
0x122: frame_vm_group_bin_6165 (RW)
0x123: frame_vm_group_bin_22347 (RW)
0x124: frame_vm_group_bin_15163 (RW)
0x125: frame_vm_group_bin_7984 (RW)
0x126: frame_vm_group_bin_0818 (RW)
0x127: frame_vm_group_bin_17013 (RW)
0x128: frame_vm_group_bin_9805 (RW)
0x129: frame_vm_group_bin_2644 (RW)
0x12: frame_vm_group_bin_21676 (RW)
0x12a: frame_vm_group_bin_18719 (RW)
0x12b: frame_vm_group_bin_11632 (RW)
0x12c: frame_vm_group_bin_4475 (RW)
0x12d: frame_vm_group_bin_20571 (RW)
0x12e: frame_vm_group_bin_9723 (RW)
0x12f: frame_vm_group_bin_6196 (RW)
0x130: frame_vm_group_bin_22380 (RW)
0x131: frame_vm_group_bin_15196 (RW)
0x132: frame_vm_group_bin_4011 (RW)
0x133: frame_vm_group_bin_0851 (RW)
0x134: frame_vm_group_bin_17046 (RW)
0x135: frame_vm_group_bin_9838 (RW)
0x136: frame_vm_group_bin_2677 (RW)
0x137: frame_vm_group_bin_18750 (RW)
0x138: frame_vm_group_bin_11655 (RW)
0x139: frame_vm_group_bin_4508 (RW)
0x13: frame_vm_group_bin_14500 (RW)
0x13a: frame_vm_group_bin_20605 (RW)
0x13b: frame_vm_group_bin_13405 (RW)
0x13c: frame_vm_group_bin_6224 (RW)
0x13d: frame_vm_group_bin_22414 (RW)
0x13e: frame_vm_group_bin_15231 (RW)
0x13f: frame_vm_group_bin_8043 (RW)
0x140: frame_vm_group_bin_0885 (RW)
0x141: frame_vm_group_bin_17080 (RW)
0x142: frame_vm_group_bin_9872 (RW)
0x143: frame_vm_group_bin_2711 (RW)
0x144: frame_vm_group_bin_18784 (RW)
0x145: frame_vm_group_bin_11679 (RW)
0x146: frame_vm_group_bin_4542 (RW)
0x147: frame_vm_group_bin_20638 (RW)
0x148: frame_vm_group_bin_13438 (RW)
0x149: frame_vm_group_bin_6254 (RW)
0x14: frame_vm_group_bin_7287 (RW)
0x14a: frame_vm_group_bin_22446 (RW)
0x14b: frame_vm_group_bin_15264 (RW)
0x14c: frame_vm_group_bin_8074 (RW)
0x14d: frame_vm_group_bin_0918 (RW)
0x14e: frame_vm_group_bin_17113 (RW)
0x14f: frame_vm_group_bin_9904 (RW)
0x150: frame_vm_group_bin_2744 (RW)
0x151: frame_vm_group_bin_18817 (RW)
0x152: frame_vm_group_bin_11706 (RW)
0x153: frame_vm_group_bin_3321 (RW)
0x154: frame_vm_group_bin_20670 (RW)
0x155: frame_vm_group_bin_13471 (RW)
0x156: frame_vm_group_bin_6286 (RW)
0x157: frame_vm_group_bin_22479 (RW)
0x158: frame_vm_group_bin_15296 (RW)
0x159: frame_vm_group_bin_8106 (RW)
0x15: frame_vm_group_bin_0163 (RW)
0x15a: frame_vm_group_bin_0952 (RW)
0x15b: frame_vm_group_bin_17147 (RW)
0x15c: frame_vm_group_bin_13664 (RW)
0x15d: frame_vm_group_bin_2778 (RW)
0x15e: frame_vm_group_bin_18852 (RW)
0x15f: frame_vm_group_bin_11732 (RW)
0x160: frame_vm_group_bin_7928 (RW)
0x161: frame_vm_group_bin_20704 (RW)
0x162: frame_vm_group_bin_13505 (RW)
0x163: frame_vm_group_bin_6319 (RW)
0x164: frame_vm_group_bin_22513 (RW)
0x165: frame_vm_group_bin_15330 (RW)
0x166: frame_vm_group_bin_8139 (RW)
0x167: frame_vm_group_bin_0985 (RW)
0x168: frame_vm_group_bin_17178 (RW)
0x169: frame_vm_group_bin_9969 (RW)
0x16: frame_vm_group_bin_16316 (RW)
0x16a: frame_vm_group_bin_2811 (RW)
0x16b: frame_vm_group_bin_18885 (RW)
0x16c: frame_vm_group_bin_11753 (RW)
0x16d: frame_vm_group_bin_4619 (RW)
0x16e: frame_vm_group_bin_20737 (RW)
0x16f: frame_vm_group_bin_13538 (RW)
0x170: frame_vm_group_bin_6352 (RW)
0x171: frame_vm_group_bin_22545 (RW)
0x172: frame_vm_group_bin_15363 (RW)
0x173: frame_vm_group_bin_8172 (RW)
0x174: frame_vm_group_bin_1017 (RW)
0x175: frame_vm_group_bin_17209 (RW)
0x176: frame_vm_group_bin_10002 (RW)
0x177: frame_vm_group_bin_2844 (RW)
0x178: frame_vm_group_bin_18918 (RW)
0x179: frame_vm_group_bin_11778 (RW)
0x17: frame_vm_group_bin_9141 (RW)
0x17a: frame_vm_group_bin_4650 (RW)
0x17b: frame_vm_group_bin_20771 (RW)
0x17c: frame_vm_group_bin_13572 (RW)
0x17d: frame_vm_group_bin_6383 (RW)
0x17e: frame_vm_group_bin_22579 (RW)
0x17f: frame_vm_group_bin_15397 (RW)
0x180: frame_vm_group_bin_8206 (RW)
0x181: frame_vm_group_bin_7197 (RW)
0x182: frame_vm_group_bin_17242 (RW)
0x183: frame_vm_group_bin_10036 (RW)
0x184: frame_vm_group_bin_2879 (RW)
0x185: frame_vm_group_bin_18951 (RW)
0x186: frame_vm_group_bin_11808 (RW)
0x187: frame_vm_group_bin_4682 (RW)
0x188: frame_vm_group_bin_20804 (RW)
0x189: frame_vm_group_bin_13605 (RW)
0x18: frame_vm_group_bin_1953 (RW)
0x18a: frame_vm_group_bin_6415 (RW)
0x18b: frame_vm_group_bin_22612 (RW)
0x18c: frame_vm_group_bin_15430 (RW)
0x18d: frame_vm_group_bin_8239 (RW)
0x18e: frame_vm_group_bin_11886 (RW)
0x18f: frame_vm_group_bin_17275 (RW)
0x190: frame_vm_group_bin_10069 (RW)
0x191: frame_vm_group_bin_2912 (RW)
0x192: frame_vm_group_bin_18982 (RW)
0x193: frame_vm_group_bin_11840 (RW)
0x194: frame_vm_group_bin_4714 (RW)
0x195: frame_vm_group_bin_20836 (RW)
0x196: frame_vm_group_bin_0412 (RW)
0x197: frame_vm_group_bin_6448 (RW)
0x198: frame_vm_group_bin_22645 (RW)
0x199: frame_vm_group_bin_15463 (RW)
0x19: frame_vm_group_bin_18051 (RW)
0x19a: frame_vm_group_bin_8272 (RW)
0x19b: frame_vm_group_bin_1088 (RW)
0x19c: frame_vm_group_bin_17309 (RW)
0x19d: frame_vm_group_bin_10103 (RW)
0x19e: frame_vm_group_bin_2946 (RW)
0x19f: frame_vm_group_bin_19016 (RW)
0x1: frame_vm_group_bin_3710 (RW)
0x1a0: frame_vm_group_bin_11870 (RW)
0x1a1: frame_vm_group_bin_4747 (RW)
0x1a2: frame_vm_group_bin_6497 (RW)
0x1a3: frame_vm_group_bin_13671 (RW)
0x1a4: frame_vm_group_bin_6482 (RW)
0x1a5: frame_vm_group_bin_22679 (RW)
0x1a6: frame_vm_group_bin_15497 (RW)
0x1a7: frame_vm_group_bin_8305 (RW)
0x1a8: frame_vm_group_bin_1116 (RW)
0x1a9: frame_vm_group_bin_17342 (RW)
0x1a: frame_vm_group_bin_10962 (RW)
0x1aa: frame_vm_group_bin_10136 (RW)
0x1ab: frame_vm_group_bin_2979 (RW)
0x1ac: frame_vm_group_bin_19049 (RW)
0x1ad: frame_vm_group_bin_11894 (RW)
0x1ae: frame_vm_group_bin_4780 (RW)
0x1af: frame_vm_group_bin_20888 (RW)
0x1b0: frame_vm_group_bin_13704 (RW)
0x1b1: frame_vm_group_bin_6515 (RW)
0x1b2: frame_vm_group_bin_22712 (RW)
0x1b3: frame_vm_group_bin_15529 (RW)
0x1b4: frame_vm_group_bin_8338 (RW)
0x1b5: frame_vm_group_bin_1149 (RW)
0x1b6: frame_vm_group_bin_17374 (RW)
0x1b7: frame_vm_group_bin_10171 (RW)
0x1b8: frame_vm_group_bin_3012 (RW)
0x1b9: frame_vm_group_bin_19082 (RW)
0x1b: frame_vm_group_bin_3777 (RW)
0x1ba: frame_vm_group_bin_11921 (RW)
0x1bb: frame_vm_group_bin_4813 (RW)
0x1bc: frame_vm_group_bin_20918 (RW)
0x1bd: frame_vm_group_bin_13737 (RW)
0x1be: frame_vm_group_bin_6549 (RW)
0x1bf: frame_vm_group_bin_22745 (RW)
0x1c0: frame_vm_group_bin_15562 (RW)
0x1c1: frame_vm_group_bin_8372 (RW)
0x1c2: frame_vm_group_bin_1183 (RW)
0x1c3: frame_vm_group_bin_5843 (RW)
0x1c4: frame_vm_group_bin_10205 (RW)
0x1c5: frame_vm_group_bin_3046 (RW)
0x1c6: frame_vm_group_bin_19115 (RW)
0x1c7: frame_vm_group_bin_11951 (RW)
0x1c8: frame_vm_group_bin_4846 (RW)
0x1c9: frame_vm_group_bin_20532 (RW)
0x1c: frame_vm_group_bin_19877 (RW)
0x1ca: frame_vm_group_bin_13771 (RW)
0x1cb: frame_vm_group_bin_6582 (RW)
0x1cc: frame_vm_group_bin_22778 (RW)
0x1cd: frame_vm_group_bin_15595 (RW)
0x1ce: frame_vm_group_bin_8405 (RW)
0x1cf: frame_vm_group_bin_1216 (RW)
0x1d0: frame_vm_group_bin_10515 (RW)
0x1d1: frame_vm_group_bin_10238 (RW)
0x1d2: frame_vm_group_bin_3079 (RW)
0x1d3: frame_vm_group_bin_19147 (RW)
0x1d4: frame_vm_group_bin_11984 (RW)
0x1d5: frame_vm_group_bin_4879 (RW)
0x1d6: frame_vm_group_bin_20972 (RW)
0x1d7: frame_vm_group_bin_13804 (RW)
0x1d8: frame_vm_group_bin_6615 (RW)
0x1d9: frame_vm_group_bin_22811 (RW)
0x1d: frame_vm_group_bin_12691 (RW)
0x1da: frame_vm_group_bin_15629 (RW)
0x1db: frame_vm_group_bin_8439 (RW)
0x1dc: frame_vm_group_bin_1249 (RW)
0x1dd: frame_vm_group_bin_17455 (RW)
0x1de: frame_vm_group_bin_10272 (RW)
0x1df: frame_vm_group_bin_12253 (RW)
0x1e0: frame_vm_group_bin_19181 (RW)
0x1e1: frame_vm_group_bin_12016 (RW)
0x1e2: frame_vm_group_bin_4913 (RW)
0x1e3: frame_vm_group_bin_21006 (RW)
0x1e4: frame_vm_group_bin_17452 (RW)
0x1e5: frame_vm_group_bin_6649 (RW)
0x1e6: frame_vm_group_bin_22845 (RW)
0x1e7: frame_vm_group_bin_15662 (RW)
0x1e8: frame_vm_group_bin_8472 (RW)
0x1e9: frame_vm_group_bin_1280 (RW)
0x1e: frame_vm_group_bin_5611 (RW)
0x1ea: frame_vm_group_bin_17473 (RW)
0x1eb: frame_vm_group_bin_10305 (RW)
0x1ec: frame_vm_group_bin_3145 (RW)
0x1ed: frame_vm_group_bin_19214 (RW)
0x1ee: frame_vm_group_bin_12046 (RW)
0x1ef: frame_vm_group_bin_4944 (RW)
0x1f0: frame_vm_group_bin_21039 (RW)
0x1f1: frame_vm_group_bin_13863 (RW)
0x1f2: frame_vm_group_bin_6682 (RW)
0x1f3: frame_vm_group_bin_22878 (RW)
0x1f4: frame_vm_group_bin_15695 (RW)
0x1f5: frame_vm_group_bin_8505 (RW)
0x1f6: frame_vm_group_bin_2631 (RW)
0x1f7: frame_vm_group_bin_17496 (RW)
0x1f8: frame_vm_group_bin_10338 (RW)
0x1f9: frame_vm_group_bin_3178 (RW)
0x1f: frame_vm_group_bin_21709 (RW)
0x1fa: frame_vm_group_bin_19248 (RW)
0x1fb: frame_vm_group_bin_12075 (RW)
0x1fc: frame_vm_group_bin_4976 (RW)
0x1fd: frame_vm_group_bin_21074 (RW)
0x1fe: frame_vm_group_bin_13896 (RW)
0x1ff: frame_vm_group_bin_6715 (RW)
0x20: frame_vm_group_bin_14535 (RW)
0x21: frame_vm_group_bin_7320 (RW)
0x22: frame_vm_group_bin_0194 (RW)
0x23: frame_vm_group_bin_16349 (RW)
0x24: frame_vm_group_bin_9173 (RW)
0x25: frame_vm_group_bin_1986 (RW)
0x26: frame_vm_group_bin_18083 (RW)
0x27: frame_vm_group_bin_10994 (RW)
0x28: frame_vm_group_bin_3809 (RW)
0x29: frame_vm_group_bin_19908 (RW)
0x2: frame_vm_group_bin_19810 (RW)
0x2a: frame_vm_group_bin_9628 (RW)
0x2b: frame_vm_group_bin_5642 (RW)
0x2c: frame_vm_group_bin_21742 (RW)
0x2d: frame_vm_group_bin_14568 (RW)
0x2e: frame_vm_group_bin_7353 (RW)
0x2f: frame_vm_group_bin_0225 (RW)
0x30: frame_vm_group_bin_16382 (RW)
0x31: frame_vm_group_bin_22931 (RW)
0x32: frame_vm_group_bin_2019 (RW)
0x33: frame_vm_group_bin_18115 (RW)
0x34: frame_vm_group_bin_11027 (RW)
0x35: frame_vm_group_bin_3842 (RW)
0x36: frame_vm_group_bin_19940 (RW)
0x37: frame_vm_group_bin_12740 (RW)
0x38: frame_vm_group_bin_5675 (RW)
0x39: frame_vm_group_bin_21775 (RW)
0x3: frame_vm_group_bin_12638 (RW)
0x3a: frame_vm_group_bin_14602 (RW)
0x3b: frame_vm_group_bin_7387 (RW)
0x3c: frame_vm_group_bin_0249 (RW)
0x3d: frame_vm_group_bin_16416 (RW)
0x3e: frame_vm_group_bin_9229 (RW)
0x3f: frame_vm_group_bin_2053 (RW)
0x40: frame_vm_group_bin_18149 (RW)
0x41: frame_vm_group_bin_11061 (RW)
0x42: frame_vm_group_bin_3876 (RW)
0x43: frame_vm_group_bin_19974 (RW)
0x44: frame_vm_group_bin_12773 (RW)
0x45: frame_vm_group_bin_5709 (RW)
0x46: frame_vm_group_bin_21809 (RW)
0x47: frame_vm_group_bin_14634 (RW)
0x48: frame_vm_group_bin_7420 (RW)
0x49: frame_vm_group_bin_0272 (RW)
0x4: frame_vm_group_bin_5545 (RW)
0x4a: frame_vm_group_bin_16449 (RW)
0x4b: frame_vm_group_bin_8929 (RW)
0x4c: frame_vm_group_bin_2086 (RW)
0x4d: frame_vm_group_bin_18182 (RW)
0x4e: frame_vm_group_bin_11094 (RW)
0x4f: frame_vm_group_bin_3909 (RW)
0x50: frame_vm_group_bin_20005 (RW)
0x51: frame_vm_group_bin_12806 (RW)
0x52: frame_vm_group_bin_5741 (RW)
0x53: frame_vm_group_bin_21842 (RW)
0x54: frame_vm_group_bin_14667 (RW)
0x55: frame_vm_group_bin_7453 (RW)
0x56: frame_vm_group_bin_0301 (RW)
0x57: frame_vm_group_bin_16482 (RW)
0x58: frame_vm_group_bin_9277 (RW)
0x59: frame_vm_group_bin_2120 (RW)
0x5: frame_vm_group_bin_21643 (RW)
0x5a: frame_vm_group_bin_18215 (RW)
0x5b: frame_vm_group_bin_11127 (RW)
0x5c: frame_vm_group_bin_3942 (RW)
0x5d: frame_vm_group_bin_20039 (RW)
0x5e: frame_vm_group_bin_12839 (RW)
0x5f: frame_vm_group_bin_5765 (RW)
0x60: frame_vm_group_bin_21876 (RW)
0x61: frame_vm_group_bin_14701 (RW)
0x62: frame_vm_group_bin_7487 (RW)
0x63: frame_vm_group_bin_0333 (RW)
0x64: frame_vm_group_bin_16516 (RW)
0x65: frame_vm_group_bin_9305 (RW)
0x66: frame_vm_group_bin_2154 (RW)
0x67: frame_vm_group_bin_18248 (RW)
0x68: frame_vm_group_bin_11160 (RW)
0x69: frame_vm_group_bin_3975 (RW)
0x6: frame_vm_group_bin_14467 (RW)
0x6a: frame_vm_group_bin_20072 (RW)
0x6b: frame_vm_group_bin_12872 (RW)
0x6c: frame_vm_group_bin_8200 (RW)
0x6d: frame_vm_group_bin_21909 (RW)
0x6e: frame_vm_group_bin_14734 (RW)
0x6f: frame_vm_group_bin_7519 (RW)
0x70: frame_vm_group_bin_0365 (RW)
0x71: frame_vm_group_bin_16549 (RW)
0x72: frame_vm_group_bin_9337 (RW)
0x73: frame_vm_group_bin_2187 (RW)
0x74: frame_vm_group_bin_18281 (RW)
0x75: frame_vm_group_bin_11193 (RW)
0x76: frame_vm_group_bin_4008 (RW)
0x77: frame_vm_group_bin_20105 (RW)
0x78: frame_vm_group_bin_12905 (RW)
0x79: frame_vm_group_bin_5809 (RW)
0x7: frame_vm_group_bin_7254 (RW)
0x7a: frame_vm_group_bin_21942 (RW)
0x7b: frame_vm_group_bin_14767 (RW)
0x7c: frame_vm_group_bin_7551 (RW)
0x7d: frame_vm_group_bin_0397 (RW)
0x7e: frame_vm_group_bin_16582 (RW)
0x7f: frame_vm_group_bin_9371 (RW)
0x80: frame_vm_group_bin_2217 (RW)
0x81: frame_vm_group_bin_18315 (RW)
0x82: frame_vm_group_bin_11227 (RW)
0x83: frame_vm_group_bin_4042 (RW)
0x84: frame_vm_group_bin_20138 (RW)
0x85: frame_vm_group_bin_12938 (RW)
0x86: frame_vm_group_bin_5834 (RW)
0x87: frame_vm_group_bin_21975 (RW)
0x88: frame_vm_group_bin_14799 (RW)
0x89: frame_vm_group_bin_7584 (RW)
0x8: frame_vm_group_bin_0141 (RW)
0x8a: frame_vm_group_bin_0424 (RW)
0x8b: frame_vm_group_bin_16614 (RW)
0x8c: frame_vm_group_bin_9405 (RW)
0x8d: frame_vm_group_bin_2245 (RW)
0x8e: frame_vm_group_bin_18348 (RW)
0x8f: frame_vm_group_bin_11260 (RW)
0x90: frame_vm_group_bin_4075 (RW)
0x91: frame_vm_group_bin_20170 (RW)
0x92: frame_vm_group_bin_12971 (RW)
0x93: frame_vm_group_bin_5858 (RW)
0x94: frame_vm_group_bin_22008 (RW)
0x95: frame_vm_group_bin_14832 (RW)
0x96: frame_vm_group_bin_7617 (RW)
0x97: frame_vm_group_bin_0457 (RW)
0x98: frame_vm_group_bin_16647 (RW)
0x99: frame_vm_group_bin_9438 (RW)
0x9: frame_vm_group_bin_16284 (RW)
0x9a: frame_vm_group_bin_2279 (RW)
0x9b: frame_vm_group_bin_18382 (RW)
0x9c: frame_vm_group_bin_11294 (RW)
0x9d: frame_vm_group_bin_4108 (RW)
0x9e: frame_vm_group_bin_20203 (RW)
0x9f: frame_vm_group_bin_13007 (RW)
0xa0: frame_vm_group_bin_5884 (RW)
0xa1: frame_vm_group_bin_2144 (RW)
0xa2: frame_vm_group_bin_14866 (RW)
0xa3: frame_vm_group_bin_7651 (RW)
0xa4: frame_vm_group_bin_0490 (RW)
0xa5: frame_vm_group_bin_16681 (RW)
0xa6: frame_vm_group_bin_9472 (RW)
0xa7: frame_vm_group_bin_2312 (RW)
0xa8: frame_vm_group_bin_18413 (RW)
0xa9: frame_vm_group_bin_11327 (RW)
0xa: frame_vm_group_bin_9108 (RW)
0xaa: frame_vm_group_bin_4141 (RW)
0xab: frame_vm_group_bin_20236 (RW)
0xac: frame_vm_group_bin_13040 (RW)
0xad: frame_vm_group_bin_5910 (RW)
0xae: frame_vm_group_bin_22055 (RW)
0xaf: frame_vm_group_bin_14899 (RW)
0xb0: frame_vm_group_bin_7684 (RW)
0xb1: frame_vm_group_bin_0523 (RW)
0xb2: frame_vm_group_bin_16713 (RW)
0xb3: frame_vm_group_bin_9505 (RW)
0xb4: frame_vm_group_bin_2345 (RW)
0xb5: frame_vm_group_bin_18446 (RW)
0xb6: frame_vm_group_bin_11358 (RW)
0xb7: frame_vm_group_bin_4173 (RW)
0xb8: frame_vm_group_bin_15794 (RW)
0xb9: frame_vm_group_bin_13073 (RW)
0xb: frame_vm_group_bin_1920 (RW)
0xba: frame_vm_group_bin_5936 (RW)
0xbb: frame_vm_group_bin_22084 (RW)
0xbc: frame_vm_group_bin_14933 (RW)
0xbd: frame_vm_group_bin_8600 (RW)
0xbe: frame_vm_group_bin_0555 (RW)
0xbf: frame_vm_group_bin_16748 (RW)
0xc0: frame_vm_group_bin_9539 (RW)
0xc1: frame_vm_group_bin_2379 (RW)
0xc2: frame_vm_group_bin_1410 (RW)
0xc3: frame_vm_group_bin_11391 (RW)
0xc4: frame_vm_group_bin_4206 (RW)
0xc5: frame_vm_group_bin_20302 (RW)
0xc6: frame_vm_group_bin_13107 (RW)
0xc7: frame_vm_group_bin_5958 (RW)
0xc8: frame_vm_group_bin_22115 (RW)
0xc9: frame_vm_group_bin_14966 (RW)
0xc: frame_vm_group_bin_18018 (RW)
0xca: frame_vm_group_bin_7750 (RW)
0xcb: frame_vm_group_bin_0586 (RW)
0xcc: frame_vm_group_bin_16781 (RW)
0xcd: frame_vm_group_bin_9572 (RW)
0xce: frame_vm_group_bin_2412 (RW)
0xcf: frame_vm_group_bin_6069 (RW)
0xd0: frame_vm_group_bin_11423 (RW)
0xd1: frame_vm_group_bin_4239 (RW)
0xd2: frame_vm_group_bin_20337 (RW)
0xd3: frame_vm_group_bin_13140 (RW)
0xd4: frame_vm_group_bin_5987 (RW)
0xd5: frame_vm_group_bin_22148 (RW)
0xd6: frame_vm_group_bin_14999 (RW)
0xd7: frame_vm_group_bin_7783 (RW)
0xd8: frame_vm_group_bin_0619 (RW)
0xd9: frame_vm_group_bin_16814 (RW)
0xd: frame_vm_group_bin_10928 (RW)
0xda: frame_vm_group_bin_9606 (RW)
0xdb: frame_vm_group_bin_2445 (RW)
0xdc: frame_vm_group_bin_18531 (RW)
0xdd: frame_vm_group_bin_11457 (RW)
0xde: frame_vm_group_bin_4273 (RW)
0xdf: frame_vm_group_bin_20371 (RW)
0xe0: frame_vm_group_bin_13174 (RW)
0xe1: frame_vm_group_bin_6018 (RW)
0xe2: frame_vm_group_bin_22182 (RW)
0xe3: frame_vm_group_bin_15033 (RW)
0xe4: frame_vm_group_bin_7817 (RW)
0xe5: frame_vm_group_bin_0652 (RW)
0xe6: frame_vm_group_bin_16848 (RW)
0xe7: frame_vm_group_bin_9639 (RW)
0xe8: frame_vm_group_bin_2477 (RW)
0xe9: frame_vm_group_bin_18556 (RW)
0xe: frame_vm_group_bin_3743 (RW)
0xea: frame_vm_group_bin_11490 (RW)
0xeb: frame_vm_group_bin_4306 (RW)
0xec: frame_vm_group_bin_20404 (RW)
0xed: frame_vm_group_bin_13207 (RW)
0xee: frame_vm_group_bin_6046 (RW)
0xef: frame_vm_group_bin_22215 (RW)
0xf0: frame_vm_group_bin_5444 (RW)
0xf1: frame_vm_group_bin_7849 (RW)
0xf2: frame_vm_group_bin_0685 (RW)
0xf3: frame_vm_group_bin_16880 (RW)
0xf4: frame_vm_group_bin_9672 (RW)
0xf5: frame_vm_group_bin_2510 (RW)
0xf6: frame_vm_group_bin_18587 (RW)
0xf7: frame_vm_group_bin_11523 (RW)
0xf8: frame_vm_group_bin_4339 (RW)
0xf9: frame_vm_group_bin_20437 (RW)
0xf: frame_vm_group_bin_19843 (RW)
0xfa: frame_vm_group_bin_13241 (RW)
0xfb: frame_vm_group_bin_6071 (RW)
0xfc: frame_vm_group_bin_22249 (RW)
0xfd: frame_vm_group_bin_15083 (RW)
0xfe: frame_vm_group_bin_7883 (RW)
0xff: frame_vm_group_bin_0719 (RW)
}
pt_vm_group_bin_0196 {
0x0: frame_vm_group_bin_14134 (RW)
0x100: frame_vm_group_bin_20134 (RW)
0x101: frame_vm_group_bin_12934 (RW)
0x102: frame_vm_group_bin_14554 (RW)
0x103: frame_vm_group_bin_21971 (RW)
0x104: frame_vm_group_bin_14795 (RW)
0x105: frame_vm_group_bin_7580 (RW)
0x106: frame_vm_group_bin_8814 (RW)
0x107: frame_vm_group_bin_16610 (RW)
0x108: frame_vm_group_bin_9401 (RW)
0x109: frame_vm_group_bin_2242 (RW)
0x10: frame_vm_group_bin_16000 (RW)
0x10a: frame_vm_group_bin_18344 (RW)
0x10b: frame_vm_group_bin_11256 (RW)
0x10c: frame_vm_group_bin_4071 (RW)
0x10d: frame_vm_group_bin_20166 (RW)
0x10e: frame_vm_group_bin_12967 (RW)
0x10f: frame_vm_group_bin_5855 (RW)
0x110: frame_vm_group_bin_22004 (RW)
0x111: frame_vm_group_bin_14828 (RW)
0x112: frame_vm_group_bin_7613 (RW)
0x113: frame_vm_group_bin_0453 (RW)
0x114: frame_vm_group_bin_16643 (RW)
0x115: frame_vm_group_bin_9434 (RW)
0x116: frame_vm_group_bin_2274 (RW)
0x117: frame_vm_group_bin_18377 (RW)
0x118: frame_vm_group_bin_11289 (RW)
0x119: frame_vm_group_bin_4104 (RW)
0x11: frame_vm_group_bin_8807 (RW)
0x11a: frame_vm_group_bin_20199 (RW)
0x11b: frame_vm_group_bin_13003 (RW)
0x11c: frame_vm_group_bin_0551 (RW)
0x11d: frame_vm_group_bin_22032 (RW)
0x11e: frame_vm_group_bin_14862 (RW)
0x11f: frame_vm_group_bin_7647 (RW)
0x120: frame_vm_group_bin_0486 (RW)
0x121: frame_vm_group_bin_16677 (RW)
0x122: frame_vm_group_bin_9468 (RW)
0x123: frame_vm_group_bin_2308 (RW)
0x124: frame_vm_group_bin_18409 (RW)
0x125: frame_vm_group_bin_11323 (RW)
0x126: frame_vm_group_bin_4137 (RW)
0x127: frame_vm_group_bin_20232 (RW)
0x128: frame_vm_group_bin_13036 (RW)
0x129: frame_vm_group_bin_5283 (RW)
0x12: frame_vm_group_bin_1618 (RW)
0x12a: frame_vm_group_bin_22053 (RW)
0x12b: frame_vm_group_bin_14895 (RW)
0x12c: frame_vm_group_bin_7680 (RW)
0x12d: frame_vm_group_bin_0519 (RW)
0x12e: frame_vm_group_bin_16709 (RW)
0x12f: frame_vm_group_bin_9501 (RW)
0x130: frame_vm_group_bin_2341 (RW)
0x131: frame_vm_group_bin_18442 (RW)
0x132: frame_vm_group_bin_11354 (RW)
0x133: frame_vm_group_bin_4169 (RW)
0x134: frame_vm_group_bin_20265 (RW)
0x135: frame_vm_group_bin_13069 (RW)
0x136: frame_vm_group_bin_9912 (RW)
0x137: frame_vm_group_bin_22079 (RW)
0x138: frame_vm_group_bin_14928 (RW)
0x139: frame_vm_group_bin_7713 (RW)
0x13: frame_vm_group_bin_7620 (RW)
0x13a: frame_vm_group_bin_4198 (RW)
0x13b: frame_vm_group_bin_16744 (RW)
0x13c: frame_vm_group_bin_9535 (RW)
0x13d: frame_vm_group_bin_2375 (RW)
0x13e: frame_vm_group_bin_18474 (RW)
0x13f: frame_vm_group_bin_11387 (RW)
0x140: frame_vm_group_bin_4202 (RW)
0x141: frame_vm_group_bin_20298 (RW)
0x142: frame_vm_group_bin_13103 (RW)
0x143: frame_vm_group_bin_14578 (RW)
0x144: frame_vm_group_bin_22111 (RW)
0x145: frame_vm_group_bin_14962 (RW)
0x146: frame_vm_group_bin_7746 (RW)
0x147: frame_vm_group_bin_8839 (RW)
0x148: frame_vm_group_bin_16777 (RW)
0x149: frame_vm_group_bin_9568 (RW)
0x14: frame_vm_group_bin_10628 (RW)
0x14a: frame_vm_group_bin_2408 (RW)
0x14b: frame_vm_group_bin_18500 (RW)
0x14c: frame_vm_group_bin_11419 (RW)
0x14d: frame_vm_group_bin_4235 (RW)
0x14e: frame_vm_group_bin_20333 (RW)
0x14f: frame_vm_group_bin_13136 (RW)
0x150: frame_vm_group_bin_5983 (RW)
0x151: frame_vm_group_bin_22144 (RW)
0x152: frame_vm_group_bin_14995 (RW)
0x153: frame_vm_group_bin_7779 (RW)
0x154: frame_vm_group_bin_0615 (RW)
0x155: frame_vm_group_bin_16810 (RW)
0x156: frame_vm_group_bin_9601 (RW)
0x157: frame_vm_group_bin_2440 (RW)
0x158: frame_vm_group_bin_18526 (RW)
0x159: frame_vm_group_bin_11452 (RW)
0x15: frame_vm_group_bin_3455 (RW)
0x15a: frame_vm_group_bin_4269 (RW)
0x15b: frame_vm_group_bin_20367 (RW)
0x15c: frame_vm_group_bin_13170 (RW)
0x15d: frame_vm_group_bin_0573 (RW)
0x15e: frame_vm_group_bin_22178 (RW)
0x15f: frame_vm_group_bin_15029 (RW)
0x160: frame_vm_group_bin_7813 (RW)
0x161: frame_vm_group_bin_0648 (RW)
0x162: frame_vm_group_bin_16844 (RW)
0x163: frame_vm_group_bin_9635 (RW)
0x164: frame_vm_group_bin_2473 (RW)
0x165: frame_vm_group_bin_18554 (RW)
0x166: frame_vm_group_bin_11486 (RW)
0x167: frame_vm_group_bin_4302 (RW)
0x168: frame_vm_group_bin_20400 (RW)
0x169: frame_vm_group_bin_13203 (RW)
0x16: frame_vm_group_bin_19548 (RW)
0x16a: frame_vm_group_bin_5306 (RW)
0x16b: frame_vm_group_bin_22211 (RW)
0x16c: frame_vm_group_bin_15054 (RW)
0x16d: frame_vm_group_bin_7845 (RW)
0x16e: frame_vm_group_bin_0681 (RW)
0x16f: frame_vm_group_bin_16876 (RW)
0x170: frame_vm_group_bin_9668 (RW)
0x171: frame_vm_group_bin_2506 (RW)
0x172: frame_vm_group_bin_18583 (RW)
0x173: frame_vm_group_bin_11519 (RW)
0x174: frame_vm_group_bin_4335 (RW)
0x175: frame_vm_group_bin_20433 (RW)
0x176: frame_vm_group_bin_13236 (RW)
0x177: frame_vm_group_bin_9935 (RW)
0x178: frame_vm_group_bin_22244 (RW)
0x179: frame_vm_group_bin_15078 (RW)
0x17: frame_vm_group_bin_12369 (RW)
0x17a: frame_vm_group_bin_7879 (RW)
0x17b: frame_vm_group_bin_0715 (RW)
0x17c: frame_vm_group_bin_16909 (RW)
0x17d: frame_vm_group_bin_9701 (RW)
0x17e: frame_vm_group_bin_2540 (RW)
0x17f: frame_vm_group_bin_18617 (RW)
0x180: frame_vm_group_bin_11553 (RW)
0x181: frame_vm_group_bin_4371 (RW)
0x182: frame_vm_group_bin_20467 (RW)
0x183: frame_vm_group_bin_13270 (RW)
0x184: frame_vm_group_bin_6097 (RW)
0x185: frame_vm_group_bin_22277 (RW)
0x186: frame_vm_group_bin_15106 (RW)
0x187: frame_vm_group_bin_7912 (RW)
0x188: frame_vm_group_bin_0748 (RW)
0x189: frame_vm_group_bin_16942 (RW)
0x18: frame_vm_group_bin_5281 (RW)
0x18a: frame_vm_group_bin_9734 (RW)
0x18b: frame_vm_group_bin_2573 (RW)
0x18c: frame_vm_group_bin_18649 (RW)
0x18d: frame_vm_group_bin_11581 (RW)
0x18e: frame_vm_group_bin_4404 (RW)
0x18f: frame_vm_group_bin_20500 (RW)
0x190: frame_vm_group_bin_13303 (RW)
0x191: frame_vm_group_bin_6128 (RW)
0x192: frame_vm_group_bin_22310 (RW)
0x193: frame_vm_group_bin_15132 (RW)
0x194: frame_vm_group_bin_7946 (RW)
0x195: frame_vm_group_bin_0781 (RW)
0x196: frame_vm_group_bin_16975 (RW)
0x197: frame_vm_group_bin_9767 (RW)
0x198: frame_vm_group_bin_2606 (RW)
0x199: frame_vm_group_bin_18682 (RW)
0x19: frame_vm_group_bin_21375 (RW)
0x19a: frame_vm_group_bin_11606 (RW)
0x19b: frame_vm_group_bin_4438 (RW)
0x19c: frame_vm_group_bin_20534 (RW)
0x19d: frame_vm_group_bin_13336 (RW)
0x19e: frame_vm_group_bin_6161 (RW)
0x19f: frame_vm_group_bin_22343 (RW)
0x1: frame_vm_group_bin_6924 (RW)
0x1a0: frame_vm_group_bin_15159 (RW)
0x1a1: frame_vm_group_bin_7980 (RW)
0x1a2: frame_vm_group_bin_0814 (RW)
0x1a3: frame_vm_group_bin_17009 (RW)
0x1a4: frame_vm_group_bin_9801 (RW)
0x1a5: frame_vm_group_bin_2640 (RW)
0x1a6: frame_vm_group_bin_18715 (RW)
0x1a7: frame_vm_group_bin_5068 (RW)
0x1a8: frame_vm_group_bin_4471 (RW)
0x1a9: frame_vm_group_bin_20567 (RW)
0x1a: frame_vm_group_bin_14200 (RW)
0x1aa: frame_vm_group_bin_13369 (RW)
0x1ab: frame_vm_group_bin_6193 (RW)
0x1ac: frame_vm_group_bin_22376 (RW)
0x1ad: frame_vm_group_bin_15192 (RW)
0x1ae: frame_vm_group_bin_8010 (RW)
0x1af: frame_vm_group_bin_0847 (RW)
0x1b0: frame_vm_group_bin_17042 (RW)
0x1b1: frame_vm_group_bin_9834 (RW)
0x1b2: frame_vm_group_bin_2673 (RW)
0x1b3: frame_vm_group_bin_18746 (RW)
0x1b4: frame_vm_group_bin_15698 (RW)
0x1b5: frame_vm_group_bin_4504 (RW)
0x1b6: frame_vm_group_bin_20600 (RW)
0x1b7: frame_vm_group_bin_13400 (RW)
0x1b8: frame_vm_group_bin_6219 (RW)
0x1b9: frame_vm_group_bin_22409 (RW)
0x1b: frame_vm_group_bin_6987 (RW)
0x1ba: frame_vm_group_bin_15227 (RW)
0x1bb: frame_vm_group_bin_8039 (RW)
0x1bc: frame_vm_group_bin_0881 (RW)
0x1bd: frame_vm_group_bin_17076 (RW)
0x1be: frame_vm_group_bin_9868 (RW)
0x1bf: frame_vm_group_bin_2707 (RW)
0x1c0: frame_vm_group_bin_18780 (RW)
0x1c1: frame_vm_group_bin_20342 (RW)
0x1c2: frame_vm_group_bin_4538 (RW)
0x1c3: frame_vm_group_bin_20634 (RW)
0x1c4: frame_vm_group_bin_13434 (RW)
0x1c5: frame_vm_group_bin_6250 (RW)
0x1c6: frame_vm_group_bin_22442 (RW)
0x1c7: frame_vm_group_bin_15260 (RW)
0x1c8: frame_vm_group_bin_8070 (RW)
0x1c9: frame_vm_group_bin_0914 (RW)
0x1c: frame_vm_group_bin_23210 (RW)
0x1ca: frame_vm_group_bin_17109 (RW)
0x1cb: frame_vm_group_bin_9900 (RW)
0x1cc: frame_vm_group_bin_2740 (RW)
0x1cd: frame_vm_group_bin_18813 (RW)
0x1ce: frame_vm_group_bin_1695 (RW)
0x1cf: frame_vm_group_bin_4569 (RW)
0x1d0: frame_vm_group_bin_20666 (RW)
0x1d1: frame_vm_group_bin_13467 (RW)
0x1d2: frame_vm_group_bin_6282 (RW)
0x1d3: frame_vm_group_bin_22475 (RW)
0x1d4: frame_vm_group_bin_15292 (RW)
0x1d5: frame_vm_group_bin_8102 (RW)
0x1d6: frame_vm_group_bin_0947 (RW)
0x1d7: frame_vm_group_bin_17142 (RW)
0x1d8: frame_vm_group_bin_9933 (RW)
0x1d9: frame_vm_group_bin_2773 (RW)
0x1d: frame_vm_group_bin_16034 (RW)
0x1da: frame_vm_group_bin_18848 (RW)
0x1db: frame_vm_group_bin_6335 (RW)
0x1dc: frame_vm_group_bin_4593 (RW)
0x1dd: frame_vm_group_bin_20700 (RW)
0x1de: frame_vm_group_bin_13501 (RW)
0x1df: frame_vm_group_bin_0621 (RW)
0x1e0: frame_vm_group_bin_22509 (RW)
0x1e1: frame_vm_group_bin_15326 (RW)
0x1e2: frame_vm_group_bin_8135 (RW)
0x1e3: frame_vm_group_bin_0981 (RW)
0x1e4: frame_vm_group_bin_17174 (RW)
0x1e5: frame_vm_group_bin_9965 (RW)
0x1e6: frame_vm_group_bin_2807 (RW)
0x1e7: frame_vm_group_bin_18881 (RW)
0x1e8: frame_vm_group_bin_11079 (RW)
0x1e9: frame_vm_group_bin_4617 (RW)
0x1e: frame_vm_group_bin_8841 (RW)
0x1ea: frame_vm_group_bin_20733 (RW)
0x1eb: frame_vm_group_bin_13534 (RW)
0x1ec: frame_vm_group_bin_6348 (RW)
0x1ed: frame_vm_group_bin_22541 (RW)
0x1ee: frame_vm_group_bin_15359 (RW)
0x1ef: frame_vm_group_bin_8168 (RW)
0x1f0: frame_vm_group_bin_1013 (RW)
0x1f1: frame_vm_group_bin_17205 (RW)
0x1f2: frame_vm_group_bin_9998 (RW)
0x1f3: frame_vm_group_bin_2840 (RW)
0x1f4: frame_vm_group_bin_18914 (RW)
0x1f5: frame_vm_group_bin_15723 (RW)
0x1f6: frame_vm_group_bin_4645 (RW)
0x1f7: frame_vm_group_bin_20766 (RW)
0x1f8: frame_vm_group_bin_13567 (RW)
0x1f9: frame_vm_group_bin_6380 (RW)
0x1f: frame_vm_group_bin_1652 (RW)
0x1fa: frame_vm_group_bin_22575 (RW)
0x1fb: frame_vm_group_bin_15393 (RW)
0x1fc: frame_vm_group_bin_8202 (RW)
0x1fd: frame_vm_group_bin_1038 (RW)
0x1fe: frame_vm_group_bin_17238 (RW)
0x1ff: frame_vm_group_bin_10032 (RW)
0x20: frame_vm_group_bin_17771 (RW)
0x21: frame_vm_group_bin_10660 (RW)
0x22: frame_vm_group_bin_3484 (RW)
0x23: frame_vm_group_bin_19583 (RW)
0x24: frame_vm_group_bin_12403 (RW)
0x25: frame_vm_group_bin_5314 (RW)
0x26: frame_vm_group_bin_21409 (RW)
0x27: frame_vm_group_bin_14233 (RW)
0x28: frame_vm_group_bin_7020 (RW)
0x29: frame_vm_group_bin_23232 (RW)
0x2: frame_vm_group_bin_23147 (RW)
0x2a: frame_vm_group_bin_16067 (RW)
0x2b: frame_vm_group_bin_8873 (RW)
0x2c: frame_vm_group_bin_1685 (RW)
0x2d: frame_vm_group_bin_17802 (RW)
0x2e: frame_vm_group_bin_10693 (RW)
0x2f: frame_vm_group_bin_3510 (RW)
0x30: frame_vm_group_bin_19616 (RW)
0x31: frame_vm_group_bin_12435 (RW)
0x32: frame_vm_group_bin_5346 (RW)
0x33: frame_vm_group_bin_21441 (RW)
0x34: frame_vm_group_bin_14265 (RW)
0x35: frame_vm_group_bin_7052 (RW)
0x36: frame_vm_group_bin_23253 (RW)
0x37: frame_vm_group_bin_16099 (RW)
0x38: frame_vm_group_bin_8905 (RW)
0x39: frame_vm_group_bin_1717 (RW)
0x3: frame_vm_group_bin_15965 (RW)
0x3a: frame_vm_group_bin_17832 (RW)
0x3b: frame_vm_group_bin_10726 (RW)
0x3c: frame_vm_group_bin_3540 (RW)
0x3d: frame_vm_group_bin_19648 (RW)
0x3e: frame_vm_group_bin_12468 (RW)
0x3f: frame_vm_group_bin_5378 (RW)
0x40: frame_vm_group_bin_21474 (RW)
0x41: frame_vm_group_bin_14297 (RW)
0x42: frame_vm_group_bin_7084 (RW)
0x43: frame_vm_group_bin_8743 (RW)
0x44: frame_vm_group_bin_16131 (RW)
0x45: frame_vm_group_bin_8938 (RW)
0x46: frame_vm_group_bin_1750 (RW)
0x47: frame_vm_group_bin_17859 (RW)
0x48: frame_vm_group_bin_10758 (RW)
0x49: frame_vm_group_bin_3571 (RW)
0x4: frame_vm_group_bin_8774 (RW)
0x4a: frame_vm_group_bin_19675 (RW)
0x4b: frame_vm_group_bin_12500 (RW)
0x4c: frame_vm_group_bin_5410 (RW)
0x4d: frame_vm_group_bin_21505 (RW)
0x4e: frame_vm_group_bin_14329 (RW)
0x4f: frame_vm_group_bin_7115 (RW)
0x50: frame_vm_group_bin_13380 (RW)
0x51: frame_vm_group_bin_16163 (RW)
0x52: frame_vm_group_bin_8970 (RW)
0x53: frame_vm_group_bin_1782 (RW)
0x54: frame_vm_group_bin_17886 (RW)
0x55: frame_vm_group_bin_10790 (RW)
0x56: frame_vm_group_bin_3605 (RW)
0x57: frame_vm_group_bin_19705 (RW)
0x58: frame_vm_group_bin_12533 (RW)
0x59: frame_vm_group_bin_5443 (RW)
0x5: frame_vm_group_bin_1585 (RW)
0x5a: frame_vm_group_bin_21539 (RW)
0x5b: frame_vm_group_bin_14363 (RW)
0x5c: frame_vm_group_bin_7148 (RW)
0x5d: frame_vm_group_bin_18029 (RW)
0x5e: frame_vm_group_bin_16197 (RW)
0x5f: frame_vm_group_bin_9004 (RW)
0x60: frame_vm_group_bin_1816 (RW)
0x61: frame_vm_group_bin_17918 (RW)
0x62: frame_vm_group_bin_10824 (RW)
0x63: frame_vm_group_bin_3639 (RW)
0x64: frame_vm_group_bin_19739 (RW)
0x65: frame_vm_group_bin_12567 (RW)
0x66: frame_vm_group_bin_5475 (RW)
0x67: frame_vm_group_bin_21572 (RW)
0x68: frame_vm_group_bin_14396 (RW)
0x69: frame_vm_group_bin_7183 (RW)
0x6: frame_vm_group_bin_3014 (RW)
0x6a: frame_vm_group_bin_22764 (RW)
0x6b: frame_vm_group_bin_16224 (RW)
0x6c: frame_vm_group_bin_9037 (RW)
0x6d: frame_vm_group_bin_1849 (RW)
0x6e: frame_vm_group_bin_17049 (RW)
0x6f: frame_vm_group_bin_10857 (RW)
0x70: frame_vm_group_bin_3672 (RW)
0x71: frame_vm_group_bin_19772 (RW)
0x72: frame_vm_group_bin_12600 (RW)
0x73: frame_vm_group_bin_5508 (RW)
0x74: frame_vm_group_bin_21605 (RW)
0x75: frame_vm_group_bin_14429 (RW)
0x76: frame_vm_group_bin_7216 (RW)
0x77: frame_vm_group_bin_4127 (RW)
0x78: frame_vm_group_bin_16250 (RW)
0x79: frame_vm_group_bin_9070 (RW)
0x7: frame_vm_group_bin_10595 (RW)
0x7a: frame_vm_group_bin_1883 (RW)
0x7b: frame_vm_group_bin_17981 (RW)
0x7c: frame_vm_group_bin_10891 (RW)
0x7d: frame_vm_group_bin_3706 (RW)
0x7e: frame_vm_group_bin_19806 (RW)
0x7f: frame_vm_group_bin_12634 (RW)
0x80: frame_vm_group_bin_5541 (RW)
0x81: frame_vm_group_bin_21639 (RW)
0x82: frame_vm_group_bin_14463 (RW)
0x83: frame_vm_group_bin_7250 (RW)
0x84: frame_vm_group_bin_8766 (RW)
0x85: frame_vm_group_bin_16281 (RW)
0x86: frame_vm_group_bin_9104 (RW)
0x87: frame_vm_group_bin_1916 (RW)
0x88: frame_vm_group_bin_18014 (RW)
0x89: frame_vm_group_bin_10924 (RW)
0x8: frame_vm_group_bin_3433 (RW)
0x8a: frame_vm_group_bin_3739 (RW)
0x8b: frame_vm_group_bin_19839 (RW)
0x8c: frame_vm_group_bin_12663 (RW)
0x8d: frame_vm_group_bin_5574 (RW)
0x8e: frame_vm_group_bin_21672 (RW)
0x8f: frame_vm_group_bin_14496 (RW)
0x90: frame_vm_group_bin_7283 (RW)
0x91: frame_vm_group_bin_0160 (RW)
0x92: frame_vm_group_bin_16312 (RW)
0x93: frame_vm_group_bin_9137 (RW)
0x94: frame_vm_group_bin_1949 (RW)
0x95: frame_vm_group_bin_18047 (RW)
0x96: frame_vm_group_bin_10957 (RW)
0x97: frame_vm_group_bin_3772 (RW)
0x98: frame_vm_group_bin_19872 (RW)
0x99: frame_vm_group_bin_12686 (RW)
0x9: frame_vm_group_bin_19515 (RW)
0x9a: frame_vm_group_bin_5607 (RW)
0x9b: frame_vm_group_bin_21705 (RW)
0x9c: frame_vm_group_bin_14531 (RW)
0x9d: frame_vm_group_bin_7316 (RW)
0x9e: frame_vm_group_bin_0191 (RW)
0x9f: frame_vm_group_bin_16345 (RW)
0xa0: frame_vm_group_bin_9169 (RW)
0xa1: frame_vm_group_bin_1982 (RW)
0xa2: frame_vm_group_bin_18079 (RW)
0xa3: frame_vm_group_bin_10990 (RW)
0xa4: frame_vm_group_bin_3805 (RW)
0xa5: frame_vm_group_bin_19904 (RW)
0xa6: frame_vm_group_bin_12714 (RW)
0xa7: frame_vm_group_bin_5638 (RW)
0xa8: frame_vm_group_bin_21738 (RW)
0xa9: frame_vm_group_bin_14564 (RW)
0xa: frame_vm_group_bin_12336 (RW)
0xaa: frame_vm_group_bin_7349 (RW)
0xab: frame_vm_group_bin_0221 (RW)
0xac: frame_vm_group_bin_16378 (RW)
0xad: frame_vm_group_bin_9200 (RW)
0xae: frame_vm_group_bin_2015 (RW)
0xaf: frame_vm_group_bin_18111 (RW)
0xb0: frame_vm_group_bin_11023 (RW)
0xb1: frame_vm_group_bin_3838 (RW)
0xb2: frame_vm_group_bin_19936 (RW)
0xb3: frame_vm_group_bin_12738 (RW)
0xb4: frame_vm_group_bin_5671 (RW)
0xb5: frame_vm_group_bin_21771 (RW)
0xb6: frame_vm_group_bin_14597 (RW)
0xb7: frame_vm_group_bin_7382 (RW)
0xb8: frame_vm_group_bin_4152 (RW)
0xb9: frame_vm_group_bin_16411 (RW)
0xb: frame_vm_group_bin_5248 (RW)
0xba: frame_vm_group_bin_9226 (RW)
0xbb: frame_vm_group_bin_2049 (RW)
0xbc: frame_vm_group_bin_18145 (RW)
0xbd: frame_vm_group_bin_11057 (RW)
0xbe: frame_vm_group_bin_3872 (RW)
0xbf: frame_vm_group_bin_19970 (RW)
0xc0: frame_vm_group_bin_12769 (RW)
0xc1: frame_vm_group_bin_5705 (RW)
0xc2: frame_vm_group_bin_21805 (RW)
0xc3: frame_vm_group_bin_14630 (RW)
0xc4: frame_vm_group_bin_7416 (RW)
0xc5: frame_vm_group_bin_0269 (RW)
0xc6: frame_vm_group_bin_16445 (RW)
0xc7: frame_vm_group_bin_9251 (RW)
0xc8: frame_vm_group_bin_2082 (RW)
0xc9: frame_vm_group_bin_18178 (RW)
0xc: frame_vm_group_bin_21342 (RW)
0xca: frame_vm_group_bin_11090 (RW)
0xcb: frame_vm_group_bin_3905 (RW)
0xcc: frame_vm_group_bin_20001 (RW)
0xcd: frame_vm_group_bin_12802 (RW)
0xce: frame_vm_group_bin_5737 (RW)
0xcf: frame_vm_group_bin_21838 (RW)
0xd0: frame_vm_group_bin_14663 (RW)
0xd1: frame_vm_group_bin_7449 (RW)
0xd2: frame_vm_group_bin_0297 (RW)
0xd3: frame_vm_group_bin_16478 (RW)
0xd4: frame_vm_group_bin_9273 (RW)
0xd5: frame_vm_group_bin_2115 (RW)
0xd6: frame_vm_group_bin_18210 (RW)
0xd7: frame_vm_group_bin_11123 (RW)
0xd8: frame_vm_group_bin_3938 (RW)
0xd9: frame_vm_group_bin_20034 (RW)
0xd: frame_vm_group_bin_14167 (RW)
0xda: frame_vm_group_bin_12835 (RW)
0xdb: frame_vm_group_bin_5763 (RW)
0xdc: frame_vm_group_bin_21872 (RW)
0xdd: frame_vm_group_bin_14697 (RW)
0xde: frame_vm_group_bin_7483 (RW)
0xdf: frame_vm_group_bin_0329 (RW)
0xe0: frame_vm_group_bin_16512 (RW)
0xe1: frame_vm_group_bin_9302 (RW)
0xe2: frame_vm_group_bin_2150 (RW)
0xe3: frame_vm_group_bin_18244 (RW)
0xe4: frame_vm_group_bin_11156 (RW)
0xe5: frame_vm_group_bin_3971 (RW)
0xe6: frame_vm_group_bin_20068 (RW)
0xe7: frame_vm_group_bin_12868 (RW)
0xe8: frame_vm_group_bin_5787 (RW)
0xe9: frame_vm_group_bin_21905 (RW)
0xe: frame_vm_group_bin_6954 (RW)
0xea: frame_vm_group_bin_14730 (RW)
0xeb: frame_vm_group_bin_7515 (RW)
0xec: frame_vm_group_bin_0361 (RW)
0xed: frame_vm_group_bin_16545 (RW)
0xee: frame_vm_group_bin_9333 (RW)
0xef: frame_vm_group_bin_2183 (RW)
0xf0: frame_vm_group_bin_18277 (RW)
0xf1: frame_vm_group_bin_11189 (RW)
0xf2: frame_vm_group_bin_4004 (RW)
0xf3: frame_vm_group_bin_20101 (RW)
0xf4: frame_vm_group_bin_12901 (RW)
0xf5: frame_vm_group_bin_9888 (RW)
0xf6: frame_vm_group_bin_21937 (RW)
0xf7: frame_vm_group_bin_14762 (RW)
0xf8: frame_vm_group_bin_7547 (RW)
0xf9: frame_vm_group_bin_0392 (RW)
0xf: frame_vm_group_bin_23180 (RW)
0xfa: frame_vm_group_bin_16578 (RW)
0xfb: frame_vm_group_bin_9367 (RW)
0xfc: frame_vm_group_bin_2213 (RW)
0xfd: frame_vm_group_bin_18311 (RW)
0xfe: frame_vm_group_bin_11223 (RW)
0xff: frame_vm_group_bin_4038 (RW)
}
pt_vm_group_bin_0203 {
0x0: frame_vm_group_bin_16346 (RW)
0x100: frame_vm_group_bin_22344 (RW)
0x101: frame_vm_group_bin_15160 (RW)
0x102: frame_vm_group_bin_7981 (RW)
0x103: frame_vm_group_bin_0815 (RW)
0x104: frame_vm_group_bin_17010 (RW)
0x105: frame_vm_group_bin_9802 (RW)
0x106: frame_vm_group_bin_2641 (RW)
0x107: frame_vm_group_bin_18716 (RW)
0x108: frame_vm_group_bin_5795 (RW)
0x109: frame_vm_group_bin_4472 (RW)
0x10: frame_vm_group_bin_18112 (RW)
0x10a: frame_vm_group_bin_20568 (RW)
0x10b: frame_vm_group_bin_13370 (RW)
0x10c: frame_vm_group_bin_0211 (RW)
0x10d: frame_vm_group_bin_22377 (RW)
0x10e: frame_vm_group_bin_15193 (RW)
0x10f: frame_vm_group_bin_8011 (RW)
0x110: frame_vm_group_bin_0848 (RW)
0x111: frame_vm_group_bin_17043 (RW)
0x112: frame_vm_group_bin_9835 (RW)
0x113: frame_vm_group_bin_2674 (RW)
0x114: frame_vm_group_bin_18747 (RW)
0x115: frame_vm_group_bin_10634 (RW)
0x116: frame_vm_group_bin_4505 (RW)
0x117: frame_vm_group_bin_20601 (RW)
0x118: frame_vm_group_bin_13401 (RW)
0x119: frame_vm_group_bin_6220 (RW)
0x11: frame_vm_group_bin_11024 (RW)
0x11a: frame_vm_group_bin_22411 (RW)
0x11b: frame_vm_group_bin_15228 (RW)
0x11c: frame_vm_group_bin_8040 (RW)
0x11d: frame_vm_group_bin_0882 (RW)
0x11e: frame_vm_group_bin_17077 (RW)
0x11f: frame_vm_group_bin_9869 (RW)
0x120: frame_vm_group_bin_2708 (RW)
0x121: frame_vm_group_bin_18781 (RW)
0x122: frame_vm_group_bin_11676 (RW)
0x123: frame_vm_group_bin_4539 (RW)
0x124: frame_vm_group_bin_20635 (RW)
0x125: frame_vm_group_bin_13435 (RW)
0x126: frame_vm_group_bin_6251 (RW)
0x127: frame_vm_group_bin_22443 (RW)
0x128: frame_vm_group_bin_15261 (RW)
0x129: frame_vm_group_bin_8071 (RW)
0x12: frame_vm_group_bin_3839 (RW)
0x12a: frame_vm_group_bin_0915 (RW)
0x12b: frame_vm_group_bin_17110 (RW)
0x12c: frame_vm_group_bin_9901 (RW)
0x12d: frame_vm_group_bin_2741 (RW)
0x12e: frame_vm_group_bin_18814 (RW)
0x12f: frame_vm_group_bin_11703 (RW)
0x130: frame_vm_group_bin_4570 (RW)
0x131: frame_vm_group_bin_20667 (RW)
0x132: frame_vm_group_bin_13468 (RW)
0x133: frame_vm_group_bin_6283 (RW)
0x134: frame_vm_group_bin_22476 (RW)
0x135: frame_vm_group_bin_15293 (RW)
0x136: frame_vm_group_bin_8103 (RW)
0x137: frame_vm_group_bin_0948 (RW)
0x138: frame_vm_group_bin_17143 (RW)
0x139: frame_vm_group_bin_9934 (RW)
0x13: frame_vm_group_bin_19937 (RW)
0x13a: frame_vm_group_bin_2775 (RW)
0x13b: frame_vm_group_bin_18849 (RW)
0x13c: frame_vm_group_bin_1269 (RW)
0x13d: frame_vm_group_bin_4594 (RW)
0x13e: frame_vm_group_bin_20701 (RW)
0x13f: frame_vm_group_bin_13502 (RW)
0x140: frame_vm_group_bin_6316 (RW)
0x141: frame_vm_group_bin_22510 (RW)
0x142: frame_vm_group_bin_15327 (RW)
0x143: frame_vm_group_bin_8136 (RW)
0x144: frame_vm_group_bin_0982 (RW)
0x145: frame_vm_group_bin_17175 (RW)
0x146: frame_vm_group_bin_9966 (RW)
0x147: frame_vm_group_bin_2808 (RW)
0x148: frame_vm_group_bin_18882 (RW)
0x149: frame_vm_group_bin_5949 (RW)
0x14: frame_vm_group_bin_12739 (RW)
0x14a: frame_vm_group_bin_4618 (RW)
0x14b: frame_vm_group_bin_20734 (RW)
0x14c: frame_vm_group_bin_13535 (RW)
0x14d: frame_vm_group_bin_6349 (RW)
0x14e: frame_vm_group_bin_22542 (RW)
0x14f: frame_vm_group_bin_15360 (RW)
0x150: frame_vm_group_bin_8169 (RW)
0x151: frame_vm_group_bin_1014 (RW)
0x152: frame_vm_group_bin_17206 (RW)
0x153: frame_vm_group_bin_9999 (RW)
0x154: frame_vm_group_bin_2841 (RW)
0x155: frame_vm_group_bin_18915 (RW)
0x156: frame_vm_group_bin_11775 (RW)
0x157: frame_vm_group_bin_4646 (RW)
0x158: frame_vm_group_bin_20767 (RW)
0x159: frame_vm_group_bin_13568 (RW)
0x15: frame_vm_group_bin_5672 (RW)
0x15a: frame_vm_group_bin_6382 (RW)
0x15b: frame_vm_group_bin_22576 (RW)
0x15c: frame_vm_group_bin_15394 (RW)
0x15d: frame_vm_group_bin_8203 (RW)
0x15e: frame_vm_group_bin_1039 (RW)
0x15f: frame_vm_group_bin_17239 (RW)
0x160: frame_vm_group_bin_10033 (RW)
0x161: frame_vm_group_bin_2876 (RW)
0x162: frame_vm_group_bin_18948 (RW)
0x163: frame_vm_group_bin_11805 (RW)
0x164: frame_vm_group_bin_4679 (RW)
0x165: frame_vm_group_bin_20801 (RW)
0x166: frame_vm_group_bin_13602 (RW)
0x167: frame_vm_group_bin_6412 (RW)
0x168: frame_vm_group_bin_22609 (RW)
0x169: frame_vm_group_bin_15427 (RW)
0x16: frame_vm_group_bin_21772 (RW)
0x16a: frame_vm_group_bin_8236 (RW)
0x16b: frame_vm_group_bin_1060 (RW)
0x16c: frame_vm_group_bin_17272 (RW)
0x16d: frame_vm_group_bin_10066 (RW)
0x16e: frame_vm_group_bin_2909 (RW)
0x16f: frame_vm_group_bin_18979 (RW)
0x170: frame_vm_group_bin_11837 (RW)
0x171: frame_vm_group_bin_4711 (RW)
0x172: frame_vm_group_bin_20833 (RW)
0x173: frame_vm_group_bin_13635 (RW)
0x174: frame_vm_group_bin_6445 (RW)
0x175: frame_vm_group_bin_22642 (RW)
0x176: frame_vm_group_bin_15460 (RW)
0x177: frame_vm_group_bin_8269 (RW)
0x178: frame_vm_group_bin_1084 (RW)
0x179: frame_vm_group_bin_17305 (RW)
0x17: frame_vm_group_bin_14598 (RW)
0x17a: frame_vm_group_bin_10100 (RW)
0x17b: frame_vm_group_bin_2943 (RW)
0x17c: frame_vm_group_bin_19013 (RW)
0x17d: frame_vm_group_bin_11867 (RW)
0x17e: frame_vm_group_bin_4744 (RW)
0x17f: frame_vm_group_bin_20862 (RW)
0x180: frame_vm_group_bin_13668 (RW)
0x181: frame_vm_group_bin_6479 (RW)
0x182: frame_vm_group_bin_22676 (RW)
0x183: frame_vm_group_bin_15494 (RW)
0x184: frame_vm_group_bin_8302 (RW)
0x185: frame_vm_group_bin_1114 (RW)
0x186: frame_vm_group_bin_17339 (RW)
0x187: frame_vm_group_bin_10133 (RW)
0x188: frame_vm_group_bin_2976 (RW)
0x189: frame_vm_group_bin_19046 (RW)
0x18: frame_vm_group_bin_7383 (RW)
0x18a: frame_vm_group_bin_5969 (RW)
0x18b: frame_vm_group_bin_4777 (RW)
0x18c: frame_vm_group_bin_20886 (RW)
0x18d: frame_vm_group_bin_13701 (RW)
0x18e: frame_vm_group_bin_6512 (RW)
0x18f: frame_vm_group_bin_22709 (RW)
0x190: frame_vm_group_bin_15526 (RW)
0x191: frame_vm_group_bin_8335 (RW)
0x192: frame_vm_group_bin_1146 (RW)
0x193: frame_vm_group_bin_17371 (RW)
0x194: frame_vm_group_bin_10168 (RW)
0x195: frame_vm_group_bin_3009 (RW)
0x196: frame_vm_group_bin_19079 (RW)
0x197: frame_vm_group_bin_10678 (RW)
0x198: frame_vm_group_bin_4810 (RW)
0x199: frame_vm_group_bin_20914 (RW)
0x19: frame_vm_group_bin_22363 (RW)
0x19a: frame_vm_group_bin_13734 (RW)
0x19b: frame_vm_group_bin_6546 (RW)
0x19c: frame_vm_group_bin_22743 (RW)
0x19d: frame_vm_group_bin_15559 (RW)
0x19e: frame_vm_group_bin_8369 (RW)
0x19f: frame_vm_group_bin_1180 (RW)
0x1: frame_vm_group_bin_9170 (RW)
0x1a0: frame_vm_group_bin_17402 (RW)
0x1a1: frame_vm_group_bin_10202 (RW)
0x1a2: frame_vm_group_bin_3043 (RW)
0x1a3: frame_vm_group_bin_19112 (RW)
0x1a4: frame_vm_group_bin_11948 (RW)
0x1a5: frame_vm_group_bin_4843 (RW)
0x1a6: frame_vm_group_bin_20944 (RW)
0x1a7: frame_vm_group_bin_13768 (RW)
0x1a8: frame_vm_group_bin_6579 (RW)
0x1a9: frame_vm_group_bin_22775 (RW)
0x1a: frame_vm_group_bin_16413 (RW)
0x1aa: frame_vm_group_bin_15592 (RW)
0x1ab: frame_vm_group_bin_8402 (RW)
0x1ac: frame_vm_group_bin_1213 (RW)
0x1ad: frame_vm_group_bin_17427 (RW)
0x1ae: frame_vm_group_bin_10235 (RW)
0x1af: frame_vm_group_bin_3076 (RW)
0x1b0: frame_vm_group_bin_19144 (RW)
0x1b1: frame_vm_group_bin_11981 (RW)
0x1b2: frame_vm_group_bin_4876 (RW)
0x1b3: frame_vm_group_bin_20969 (RW)
0x1b4: frame_vm_group_bin_13801 (RW)
0x1b5: frame_vm_group_bin_6612 (RW)
0x1b6: frame_vm_group_bin_22808 (RW)
0x1b7: frame_vm_group_bin_15625 (RW)
0x1b8: frame_vm_group_bin_8435 (RW)
0x1b9: frame_vm_group_bin_1246 (RW)
0x1b: frame_vm_group_bin_9227 (RW)
0x1ba: frame_vm_group_bin_18822 (RW)
0x1bb: frame_vm_group_bin_10269 (RW)
0x1bc: frame_vm_group_bin_3110 (RW)
0x1bd: frame_vm_group_bin_19178 (RW)
0x1be: frame_vm_group_bin_1315 (RW)
0x1bf: frame_vm_group_bin_4910 (RW)
0x1c0: frame_vm_group_bin_21003 (RW)
0x1c1: frame_vm_group_bin_13833 (RW)
0x1c2: frame_vm_group_bin_6646 (RW)
0x1c3: frame_vm_group_bin_22842 (RW)
0x1c4: frame_vm_group_bin_15659 (RW)
0x1c5: frame_vm_group_bin_8469 (RW)
0x1c6: frame_vm_group_bin_1277 (RW)
0x1c7: frame_vm_group_bin_11746 (RW)
0x1c8: frame_vm_group_bin_10302 (RW)
0x1c9: frame_vm_group_bin_3142 (RW)
0x1c: frame_vm_group_bin_2050 (RW)
0x1ca: frame_vm_group_bin_19211 (RW)
0x1cb: frame_vm_group_bin_12043 (RW)
0x1cc: frame_vm_group_bin_4941 (RW)
0x1cd: frame_vm_group_bin_21036 (RW)
0x1ce: frame_vm_group_bin_13862 (RW)
0x1cf: frame_vm_group_bin_6679 (RW)
0x1d0: frame_vm_group_bin_22875 (RW)
0x1d1: frame_vm_group_bin_15692 (RW)
0x1d2: frame_vm_group_bin_8502 (RW)
0x1d3: frame_vm_group_bin_1310 (RW)
0x1d4: frame_vm_group_bin_16435 (RW)
0x1d5: frame_vm_group_bin_10335 (RW)
0x1d6: frame_vm_group_bin_3175 (RW)
0x1d7: frame_vm_group_bin_19244 (RW)
0x1d8: frame_vm_group_bin_12071 (RW)
0x1d9: frame_vm_group_bin_4972 (RW)
0x1d: frame_vm_group_bin_18146 (RW)
0x1da: frame_vm_group_bin_21071 (RW)
0x1db: frame_vm_group_bin_13893 (RW)
0x1dc: frame_vm_group_bin_6713 (RW)
0x1dd: frame_vm_group_bin_22909 (RW)
0x1de: frame_vm_group_bin_15726 (RW)
0x1df: frame_vm_group_bin_8535 (RW)
0x1e0: frame_vm_group_bin_1343 (RW)
0x1e1: frame_vm_group_bin_21070 (RW)
0x1e2: frame_vm_group_bin_10369 (RW)
0x1e3: frame_vm_group_bin_3209 (RW)
0x1e4: frame_vm_group_bin_19278 (RW)
0x1e5: frame_vm_group_bin_12105 (RW)
0x1e6: frame_vm_group_bin_5006 (RW)
0x1e7: frame_vm_group_bin_21104 (RW)
0x1e8: frame_vm_group_bin_13926 (RW)
0x1e9: frame_vm_group_bin_6745 (RW)
0x1e: frame_vm_group_bin_11058 (RW)
0x1ea: frame_vm_group_bin_22942 (RW)
0x1eb: frame_vm_group_bin_15759 (RW)
0x1ec: frame_vm_group_bin_8566 (RW)
0x1ed: frame_vm_group_bin_1377 (RW)
0x1ee: frame_vm_group_bin_2443 (RW)
0x1ef: frame_vm_group_bin_10398 (RW)
0x1f0: frame_vm_group_bin_3241 (RW)
0x1f1: frame_vm_group_bin_19311 (RW)
0x1f2: frame_vm_group_bin_12137 (RW)
0x1f3: frame_vm_group_bin_5039 (RW)
0x1f4: frame_vm_group_bin_21137 (RW)
0x1f5: frame_vm_group_bin_13959 (RW)
0x1f6: frame_vm_group_bin_6777 (RW)
0x1f7: frame_vm_group_bin_22974 (RW)
0x1f8: frame_vm_group_bin_15792 (RW)
0x1f9: frame_vm_group_bin_8599 (RW)
0x1f: frame_vm_group_bin_3873 (RW)
0x1fa: frame_vm_group_bin_1411 (RW)
0x1fb: frame_vm_group_bin_7056 (RW)
0x1fc: frame_vm_group_bin_10425 (RW)
0x1fd: frame_vm_group_bin_3275 (RW)
0x1fe: frame_vm_group_bin_19345 (RW)
0x1ff: frame_vm_group_bin_12168 (RW)
0x20: frame_vm_group_bin_19971 (RW)
0x21: frame_vm_group_bin_12770 (RW)
0x22: frame_vm_group_bin_5706 (RW)
0x23: frame_vm_group_bin_21806 (RW)
0x24: frame_vm_group_bin_14631 (RW)
0x25: frame_vm_group_bin_7417 (RW)
0x26: frame_vm_group_bin_3728 (RW)
0x27: frame_vm_group_bin_16446 (RW)
0x28: frame_vm_group_bin_9252 (RW)
0x29: frame_vm_group_bin_2083 (RW)
0x2: frame_vm_group_bin_1983 (RW)
0x2a: frame_vm_group_bin_18179 (RW)
0x2b: frame_vm_group_bin_11091 (RW)
0x2c: frame_vm_group_bin_3906 (RW)
0x2d: frame_vm_group_bin_20002 (RW)
0x2e: frame_vm_group_bin_12803 (RW)
0x2f: frame_vm_group_bin_5738 (RW)
0x30: frame_vm_group_bin_21839 (RW)
0x31: frame_vm_group_bin_14664 (RW)
0x32: frame_vm_group_bin_7450 (RW)
0x33: frame_vm_group_bin_0298 (RW)
0x34: frame_vm_group_bin_16479 (RW)
0x35: frame_vm_group_bin_9274 (RW)
0x36: frame_vm_group_bin_2116 (RW)
0x37: frame_vm_group_bin_18211 (RW)
0x38: frame_vm_group_bin_11124 (RW)
0x39: frame_vm_group_bin_3939 (RW)
0x3: frame_vm_group_bin_18080 (RW)
0x3a: frame_vm_group_bin_20036 (RW)
0x3b: frame_vm_group_bin_12836 (RW)
0x3c: frame_vm_group_bin_5764 (RW)
0x3d: frame_vm_group_bin_21873 (RW)
0x3e: frame_vm_group_bin_14698 (RW)
0x3f: frame_vm_group_bin_7484 (RW)
0x40: frame_vm_group_bin_0330 (RW)
0x41: frame_vm_group_bin_16513 (RW)
0x42: frame_vm_group_bin_9303 (RW)
0x43: frame_vm_group_bin_2151 (RW)
0x44: frame_vm_group_bin_18245 (RW)
0x45: frame_vm_group_bin_11157 (RW)
0x46: frame_vm_group_bin_3972 (RW)
0x47: frame_vm_group_bin_20069 (RW)
0x48: frame_vm_group_bin_12869 (RW)
0x49: frame_vm_group_bin_5788 (RW)
0x4: frame_vm_group_bin_10991 (RW)
0x4a: frame_vm_group_bin_21906 (RW)
0x4b: frame_vm_group_bin_14731 (RW)
0x4c: frame_vm_group_bin_7516 (RW)
0x4d: frame_vm_group_bin_0362 (RW)
0x4e: frame_vm_group_bin_16546 (RW)
0x4f: frame_vm_group_bin_9334 (RW)
0x50: frame_vm_group_bin_2184 (RW)
0x51: frame_vm_group_bin_18278 (RW)
0x52: frame_vm_group_bin_11190 (RW)
0x53: frame_vm_group_bin_4005 (RW)
0x54: frame_vm_group_bin_20102 (RW)
0x55: frame_vm_group_bin_12902 (RW)
0x56: frame_vm_group_bin_15980 (RW)
0x57: frame_vm_group_bin_21938 (RW)
0x58: frame_vm_group_bin_14763 (RW)
0x59: frame_vm_group_bin_7548 (RW)
0x5: frame_vm_group_bin_3806 (RW)
0x5a: frame_vm_group_bin_0394 (RW)
0x5b: frame_vm_group_bin_16579 (RW)
0x5c: frame_vm_group_bin_9368 (RW)
0x5d: frame_vm_group_bin_2214 (RW)
0x5e: frame_vm_group_bin_18312 (RW)
0x5f: frame_vm_group_bin_11224 (RW)
0x60: frame_vm_group_bin_4039 (RW)
0x61: frame_vm_group_bin_20135 (RW)
0x62: frame_vm_group_bin_12935 (RW)
0x63: frame_vm_group_bin_9462 (RW)
0x64: frame_vm_group_bin_21972 (RW)
0x65: frame_vm_group_bin_14796 (RW)
0x66: frame_vm_group_bin_7581 (RW)
0x67: frame_vm_group_bin_0421 (RW)
0x68: frame_vm_group_bin_16611 (RW)
0x69: frame_vm_group_bin_9402 (RW)
0x6: frame_vm_group_bin_19905 (RW)
0x6a: frame_vm_group_bin_2243 (RW)
0x6b: frame_vm_group_bin_18345 (RW)
0x6c: frame_vm_group_bin_11257 (RW)
0x6d: frame_vm_group_bin_4072 (RW)
0x6e: frame_vm_group_bin_20167 (RW)
0x6f: frame_vm_group_bin_12968 (RW)
0x70: frame_vm_group_bin_14130 (RW)
0x71: frame_vm_group_bin_22005 (RW)
0x72: frame_vm_group_bin_14829 (RW)
0x73: frame_vm_group_bin_7614 (RW)
0x74: frame_vm_group_bin_0454 (RW)
0x75: frame_vm_group_bin_16644 (RW)
0x76: frame_vm_group_bin_9435 (RW)
0x77: frame_vm_group_bin_2275 (RW)
0x78: frame_vm_group_bin_18378 (RW)
0x79: frame_vm_group_bin_11290 (RW)
0x7: frame_vm_group_bin_12715 (RW)
0x7a: frame_vm_group_bin_4106 (RW)
0x7b: frame_vm_group_bin_20200 (RW)
0x7c: frame_vm_group_bin_13004 (RW)
0x7d: frame_vm_group_bin_18753 (RW)
0x7e: frame_vm_group_bin_22033 (RW)
0x7f: frame_vm_group_bin_14863 (RW)
0x80: frame_vm_group_bin_7648 (RW)
0x81: frame_vm_group_bin_0487 (RW)
0x82: frame_vm_group_bin_16678 (RW)
0x83: frame_vm_group_bin_9469 (RW)
0x84: frame_vm_group_bin_2309 (RW)
0x85: frame_vm_group_bin_18410 (RW)
0x86: frame_vm_group_bin_11324 (RW)
0x87: frame_vm_group_bin_4138 (RW)
0x88: frame_vm_group_bin_20233 (RW)
0x89: frame_vm_group_bin_13037 (RW)
0x8: frame_vm_group_bin_5639 (RW)
0x8a: frame_vm_group_bin_0166 (RW)
0x8b: frame_vm_group_bin_22054 (RW)
0x8c: frame_vm_group_bin_14896 (RW)
0x8d: frame_vm_group_bin_7681 (RW)
0x8e: frame_vm_group_bin_0520 (RW)
0x8f: frame_vm_group_bin_16710 (RW)
0x90: frame_vm_group_bin_9502 (RW)
0x91: frame_vm_group_bin_2342 (RW)
0x92: frame_vm_group_bin_18443 (RW)
0x93: frame_vm_group_bin_11355 (RW)
0x94: frame_vm_group_bin_4170 (RW)
0x95: frame_vm_group_bin_20266 (RW)
0x96: frame_vm_group_bin_13070 (RW)
0x97: frame_vm_group_bin_4857 (RW)
0x98: frame_vm_group_bin_22080 (RW)
0x99: frame_vm_group_bin_14929 (RW)
0x9: frame_vm_group_bin_21739 (RW)
0x9a: frame_vm_group_bin_7715 (RW)
0x9b: frame_vm_group_bin_0552 (RW)
0x9c: frame_vm_group_bin_16745 (RW)
0x9d: frame_vm_group_bin_9536 (RW)
0x9e: frame_vm_group_bin_2376 (RW)
0x9f: frame_vm_group_bin_18475 (RW)
0xa0: frame_vm_group_bin_11388 (RW)
0xa1: frame_vm_group_bin_4203 (RW)
0xa2: frame_vm_group_bin_20299 (RW)
0xa3: frame_vm_group_bin_13104 (RW)
0xa4: frame_vm_group_bin_5955 (RW)
0xa5: frame_vm_group_bin_22112 (RW)
0xa6: frame_vm_group_bin_14963 (RW)
0xa7: frame_vm_group_bin_7747 (RW)
0xa8: frame_vm_group_bin_0583 (RW)
0xa9: frame_vm_group_bin_16778 (RW)
0xa: frame_vm_group_bin_14565 (RW)
0xaa: frame_vm_group_bin_9569 (RW)
0xab: frame_vm_group_bin_2409 (RW)
0xac: frame_vm_group_bin_18501 (RW)
0xad: frame_vm_group_bin_11420 (RW)
0xae: frame_vm_group_bin_4236 (RW)
0xaf: frame_vm_group_bin_20334 (RW)
0xb0: frame_vm_group_bin_13137 (RW)
0xb1: frame_vm_group_bin_5984 (RW)
0xb2: frame_vm_group_bin_22145 (RW)
0xb3: frame_vm_group_bin_14996 (RW)
0xb4: frame_vm_group_bin_7780 (RW)
0xb5: frame_vm_group_bin_0616 (RW)
0xb6: frame_vm_group_bin_16811 (RW)
0xb7: frame_vm_group_bin_9602 (RW)
0xb8: frame_vm_group_bin_2441 (RW)
0xb9: frame_vm_group_bin_18527 (RW)
0xb: frame_vm_group_bin_7350 (RW)
0xba: frame_vm_group_bin_11454 (RW)
0xbb: frame_vm_group_bin_4270 (RW)
0xbc: frame_vm_group_bin_20368 (RW)
0xbd: frame_vm_group_bin_13171 (RW)
0xbe: frame_vm_group_bin_6015 (RW)
0xbf: frame_vm_group_bin_22179 (RW)
0xc0: frame_vm_group_bin_15030 (RW)
0xc1: frame_vm_group_bin_7814 (RW)
0xc2: frame_vm_group_bin_0649 (RW)
0xc3: frame_vm_group_bin_16845 (RW)
0xc4: frame_vm_group_bin_9636 (RW)
0xc5: frame_vm_group_bin_2474 (RW)
0xc6: frame_vm_group_bin_18555 (RW)
0xc7: frame_vm_group_bin_11487 (RW)
0xc8: frame_vm_group_bin_4303 (RW)
0xc9: frame_vm_group_bin_20401 (RW)
0xc: frame_vm_group_bin_0222 (RW)
0xca: frame_vm_group_bin_13204 (RW)
0xcb: frame_vm_group_bin_0189 (RW)
0xcc: frame_vm_group_bin_22212 (RW)
0xcd: frame_vm_group_bin_15055 (RW)
0xce: frame_vm_group_bin_7846 (RW)
0xcf: frame_vm_group_bin_0682 (RW)
0xd0: frame_vm_group_bin_16877 (RW)
0xd1: frame_vm_group_bin_9669 (RW)
0xd2: frame_vm_group_bin_2507 (RW)
0xd3: frame_vm_group_bin_18584 (RW)
0xd4: frame_vm_group_bin_11520 (RW)
0xd5: frame_vm_group_bin_4336 (RW)
0xd6: frame_vm_group_bin_20434 (RW)
0xd7: frame_vm_group_bin_13237 (RW)
0xd8: frame_vm_group_bin_6067 (RW)
0xd9: frame_vm_group_bin_22245 (RW)
0xd: frame_vm_group_bin_16379 (RW)
0xda: frame_vm_group_bin_15080 (RW)
0xdb: frame_vm_group_bin_7880 (RW)
0xdc: frame_vm_group_bin_0716 (RW)
0xdd: frame_vm_group_bin_16910 (RW)
0xde: frame_vm_group_bin_9702 (RW)
0xdf: frame_vm_group_bin_2541 (RW)
0xe0: frame_vm_group_bin_18618 (RW)
0xe1: frame_vm_group_bin_11554 (RW)
0xe2: frame_vm_group_bin_4372 (RW)
0xe3: frame_vm_group_bin_20468 (RW)
0xe4: frame_vm_group_bin_13271 (RW)
0xe5: frame_vm_group_bin_6098 (RW)
0xe6: frame_vm_group_bin_22278 (RW)
0xe7: frame_vm_group_bin_15107 (RW)
0xe8: frame_vm_group_bin_7913 (RW)
0xe9: frame_vm_group_bin_0749 (RW)
0xe: frame_vm_group_bin_9201 (RW)
0xea: frame_vm_group_bin_16943 (RW)
0xeb: frame_vm_group_bin_9735 (RW)
0xec: frame_vm_group_bin_2574 (RW)
0xed: frame_vm_group_bin_18650 (RW)
0xee: frame_vm_group_bin_11582 (RW)
0xef: frame_vm_group_bin_4405 (RW)
0xf0: frame_vm_group_bin_20501 (RW)
0xf1: frame_vm_group_bin_13304 (RW)
0xf2: frame_vm_group_bin_6129 (RW)
0xf3: frame_vm_group_bin_22311 (RW)
0xf4: frame_vm_group_bin_15133 (RW)
0xf5: frame_vm_group_bin_7947 (RW)
0xf6: frame_vm_group_bin_0782 (RW)
0xf7: frame_vm_group_bin_16976 (RW)
0xf8: frame_vm_group_bin_9768 (RW)
0xf9: frame_vm_group_bin_2607 (RW)
0xf: frame_vm_group_bin_2016 (RW)
0xfa: frame_vm_group_bin_18684 (RW)
0xfb: frame_vm_group_bin_11607 (RW)
0xfc: frame_vm_group_bin_4439 (RW)
0xfd: frame_vm_group_bin_20535 (RW)
0xfe: frame_vm_group_bin_13337 (RW)
0xff: frame_vm_group_bin_6162 (RW)
}
pt_vm_group_bin_0210 {
0x0: frame_vm_group_bin_14512 (RW)
0x100: frame_vm_group_bin_20515 (RW)
0x101: frame_vm_group_bin_13317 (RW)
0x102: frame_vm_group_bin_6142 (RW)
0x103: frame_vm_group_bin_22325 (RW)
0x104: frame_vm_group_bin_15141 (RW)
0x105: frame_vm_group_bin_7961 (RW)
0x106: frame_vm_group_bin_0796 (RW)
0x107: frame_vm_group_bin_16990 (RW)
0x108: frame_vm_group_bin_9782 (RW)
0x109: frame_vm_group_bin_2621 (RW)
0x10: frame_vm_group_bin_16359 (RW)
0x10a: frame_vm_group_bin_18697 (RW)
0x10b: frame_vm_group_bin_11618 (RW)
0x10c: frame_vm_group_bin_4452 (RW)
0x10d: frame_vm_group_bin_20548 (RW)
0x10e: frame_vm_group_bin_13350 (RW)
0x10f: frame_vm_group_bin_6175 (RW)
0x110: frame_vm_group_bin_22357 (RW)
0x111: frame_vm_group_bin_15173 (RW)
0x112: frame_vm_group_bin_3297 (RW)
0x113: frame_vm_group_bin_0828 (RW)
0x114: frame_vm_group_bin_17023 (RW)
0x115: frame_vm_group_bin_9815 (RW)
0x116: frame_vm_group_bin_2654 (RW)
0x117: frame_vm_group_bin_18729 (RW)
0x118: frame_vm_group_bin_11639 (RW)
0x119: frame_vm_group_bin_4485 (RW)
0x11: frame_vm_group_bin_4341 (RW)
0x11a: frame_vm_group_bin_20582 (RW)
0x11b: frame_vm_group_bin_13382 (RW)
0x11c: frame_vm_group_bin_6206 (RW)
0x11d: frame_vm_group_bin_22391 (RW)
0x11e: frame_vm_group_bin_15207 (RW)
0x11f: frame_vm_group_bin_8024 (RW)
0x120: frame_vm_group_bin_0862 (RW)
0x121: frame_vm_group_bin_17057 (RW)
0x122: frame_vm_group_bin_9849 (RW)
0x123: frame_vm_group_bin_2688 (RW)
0x124: frame_vm_group_bin_18761 (RW)
0x125: frame_vm_group_bin_11663 (RW)
0x126: frame_vm_group_bin_4519 (RW)
0x127: frame_vm_group_bin_20615 (RW)
0x128: frame_vm_group_bin_13415 (RW)
0x129: frame_vm_group_bin_6233 (RW)
0x12: frame_vm_group_bin_1996 (RW)
0x12a: frame_vm_group_bin_22423 (RW)
0x12b: frame_vm_group_bin_15241 (RW)
0x12c: frame_vm_group_bin_8052 (RW)
0x12d: frame_vm_group_bin_0895 (RW)
0x12e: frame_vm_group_bin_17090 (RW)
0x12f: frame_vm_group_bin_9882 (RW)
0x130: frame_vm_group_bin_2721 (RW)
0x131: frame_vm_group_bin_18794 (RW)
0x132: frame_vm_group_bin_11687 (RW)
0x133: frame_vm_group_bin_13756 (RW)
0x134: frame_vm_group_bin_20648 (RW)
0x135: frame_vm_group_bin_13448 (RW)
0x136: frame_vm_group_bin_6264 (RW)
0x137: frame_vm_group_bin_22456 (RW)
0x138: frame_vm_group_bin_15274 (RW)
0x139: frame_vm_group_bin_8083 (RW)
0x13: frame_vm_group_bin_18093 (RW)
0x13a: frame_vm_group_bin_0929 (RW)
0x13b: frame_vm_group_bin_17124 (RW)
0x13c: frame_vm_group_bin_9915 (RW)
0x13d: frame_vm_group_bin_2755 (RW)
0x13e: frame_vm_group_bin_18829 (RW)
0x13f: frame_vm_group_bin_11716 (RW)
0x140: frame_vm_group_bin_7173 (RW)
0x141: frame_vm_group_bin_20681 (RW)
0x142: frame_vm_group_bin_13482 (RW)
0x143: frame_vm_group_bin_6297 (RW)
0x144: frame_vm_group_bin_22490 (RW)
0x145: frame_vm_group_bin_15307 (RW)
0x146: frame_vm_group_bin_8116 (RW)
0x147: frame_vm_group_bin_0962 (RW)
0x148: frame_vm_group_bin_17156 (RW)
0x149: frame_vm_group_bin_9946 (RW)
0x14: frame_vm_group_bin_11004 (RW)
0x14a: frame_vm_group_bin_2788 (RW)
0x14b: frame_vm_group_bin_18862 (RW)
0x14c: frame_vm_group_bin_11740 (RW)
0x14d: frame_vm_group_bin_4602 (RW)
0x14e: frame_vm_group_bin_20714 (RW)
0x14f: frame_vm_group_bin_13515 (RW)
0x150: frame_vm_group_bin_6329 (RW)
0x151: frame_vm_group_bin_22523 (RW)
0x152: frame_vm_group_bin_15340 (RW)
0x153: frame_vm_group_bin_8149 (RW)
0x154: frame_vm_group_bin_0995 (RW)
0x155: frame_vm_group_bin_17188 (RW)
0x156: frame_vm_group_bin_9979 (RW)
0x157: frame_vm_group_bin_2821 (RW)
0x158: frame_vm_group_bin_18895 (RW)
0x159: frame_vm_group_bin_11761 (RW)
0x15: frame_vm_group_bin_3819 (RW)
0x15a: frame_vm_group_bin_4628 (RW)
0x15b: frame_vm_group_bin_20748 (RW)
0x15c: frame_vm_group_bin_13549 (RW)
0x15d: frame_vm_group_bin_6363 (RW)
0x15e: frame_vm_group_bin_22556 (RW)
0x15f: frame_vm_group_bin_15374 (RW)
0x160: frame_vm_group_bin_8183 (RW)
0x161: frame_vm_group_bin_6474 (RW)
0x162: frame_vm_group_bin_17220 (RW)
0x163: frame_vm_group_bin_10013 (RW)
0x164: frame_vm_group_bin_2855 (RW)
0x165: frame_vm_group_bin_18929 (RW)
0x166: frame_vm_group_bin_11787 (RW)
0x167: frame_vm_group_bin_4660 (RW)
0x168: frame_vm_group_bin_20781 (RW)
0x169: frame_vm_group_bin_13582 (RW)
0x16: frame_vm_group_bin_19918 (RW)
0x16a: frame_vm_group_bin_6393 (RW)
0x16b: frame_vm_group_bin_22589 (RW)
0x16c: frame_vm_group_bin_15407 (RW)
0x16d: frame_vm_group_bin_8216 (RW)
0x16e: frame_vm_group_bin_11221 (RW)
0x16f: frame_vm_group_bin_17252 (RW)
0x170: frame_vm_group_bin_10046 (RW)
0x171: frame_vm_group_bin_2889 (RW)
0x172: frame_vm_group_bin_18961 (RW)
0x173: frame_vm_group_bin_11818 (RW)
0x174: frame_vm_group_bin_4692 (RW)
0x175: frame_vm_group_bin_20814 (RW)
0x176: frame_vm_group_bin_13615 (RW)
0x177: frame_vm_group_bin_6425 (RW)
0x178: frame_vm_group_bin_22622 (RW)
0x179: frame_vm_group_bin_15440 (RW)
0x17: frame_vm_group_bin_12722 (RW)
0x17a: frame_vm_group_bin_8250 (RW)
0x17b: frame_vm_group_bin_1070 (RW)
0x17c: frame_vm_group_bin_17286 (RW)
0x17d: frame_vm_group_bin_10080 (RW)
0x17e: frame_vm_group_bin_2923 (RW)
0x17f: frame_vm_group_bin_18993 (RW)
0x180: frame_vm_group_bin_11849 (RW)
0x181: frame_vm_group_bin_4724 (RW)
0x182: frame_vm_group_bin_5826 (RW)
0x183: frame_vm_group_bin_13648 (RW)
0x184: frame_vm_group_bin_6459 (RW)
0x185: frame_vm_group_bin_22656 (RW)
0x186: frame_vm_group_bin_15474 (RW)
0x187: frame_vm_group_bin_8282 (RW)
0x188: frame_vm_group_bin_1096 (RW)
0x189: frame_vm_group_bin_17319 (RW)
0x18: frame_vm_group_bin_5652 (RW)
0x18a: frame_vm_group_bin_10113 (RW)
0x18b: frame_vm_group_bin_2956 (RW)
0x18c: frame_vm_group_bin_19026 (RW)
0x18d: frame_vm_group_bin_11878 (RW)
0x18e: frame_vm_group_bin_4757 (RW)
0x18f: frame_vm_group_bin_20869 (RW)
0x190: frame_vm_group_bin_13681 (RW)
0x191: frame_vm_group_bin_6492 (RW)
0x192: frame_vm_group_bin_22689 (RW)
0x193: frame_vm_group_bin_15507 (RW)
0x194: frame_vm_group_bin_8315 (RW)
0x195: frame_vm_group_bin_1126 (RW)
0x196: frame_vm_group_bin_17352 (RW)
0x197: frame_vm_group_bin_10146 (RW)
0x198: frame_vm_group_bin_2989 (RW)
0x199: frame_vm_group_bin_19059 (RW)
0x19: frame_vm_group_bin_21752 (RW)
0x19a: frame_vm_group_bin_11902 (RW)
0x19b: frame_vm_group_bin_4791 (RW)
0x19c: frame_vm_group_bin_20899 (RW)
0x19d: frame_vm_group_bin_13714 (RW)
0x19e: frame_vm_group_bin_6526 (RW)
0x19f: frame_vm_group_bin_22723 (RW)
0x1: frame_vm_group_bin_7297 (RW)
0x1a0: frame_vm_group_bin_15539 (RW)
0x1a1: frame_vm_group_bin_8349 (RW)
0x1a2: frame_vm_group_bin_1160 (RW)
0x1a3: frame_vm_group_bin_5140 (RW)
0x1a4: frame_vm_group_bin_10182 (RW)
0x1a5: frame_vm_group_bin_3023 (RW)
0x1a6: frame_vm_group_bin_19093 (RW)
0x1a7: frame_vm_group_bin_11931 (RW)
0x1a8: frame_vm_group_bin_4823 (RW)
0x1a9: frame_vm_group_bin_20924 (RW)
0x1a: frame_vm_group_bin_14579 (RW)
0x1aa: frame_vm_group_bin_13747 (RW)
0x1ab: frame_vm_group_bin_6559 (RW)
0x1ac: frame_vm_group_bin_22755 (RW)
0x1ad: frame_vm_group_bin_15572 (RW)
0x1ae: frame_vm_group_bin_8382 (RW)
0x1af: frame_vm_group_bin_1193 (RW)
0x1b0: frame_vm_group_bin_17410 (RW)
0x1b1: frame_vm_group_bin_10215 (RW)
0x1b2: frame_vm_group_bin_3056 (RW)
0x1b3: frame_vm_group_bin_19125 (RW)
0x1b4: frame_vm_group_bin_11961 (RW)
0x1b5: frame_vm_group_bin_4856 (RW)
0x1b6: frame_vm_group_bin_20951 (RW)
0x1b7: frame_vm_group_bin_13781 (RW)
0x1b8: frame_vm_group_bin_6592 (RW)
0x1b9: frame_vm_group_bin_22788 (RW)
0x1b: frame_vm_group_bin_7364 (RW)
0x1ba: frame_vm_group_bin_15606 (RW)
0x1bb: frame_vm_group_bin_8416 (RW)
0x1bc: frame_vm_group_bin_1227 (RW)
0x1bd: frame_vm_group_bin_17438 (RW)
0x1be: frame_vm_group_bin_10249 (RW)
0x1bf: frame_vm_group_bin_3090 (RW)
0x1c0: frame_vm_group_bin_19158 (RW)
0x1c1: frame_vm_group_bin_11994 (RW)
0x1c2: frame_vm_group_bin_4890 (RW)
0x1c3: frame_vm_group_bin_20983 (RW)
0x1c4: frame_vm_group_bin_2868 (RW)
0x1c5: frame_vm_group_bin_6626 (RW)
0x1c6: frame_vm_group_bin_22822 (RW)
0x1c7: frame_vm_group_bin_15639 (RW)
0x1c8: frame_vm_group_bin_8449 (RW)
0x1c9: frame_vm_group_bin_1259 (RW)
0x1c: frame_vm_group_bin_0234 (RW)
0x1ca: frame_vm_group_bin_17460 (RW)
0x1cb: frame_vm_group_bin_10282 (RW)
0x1cc: frame_vm_group_bin_3122 (RW)
0x1cd: frame_vm_group_bin_19191 (RW)
0x1ce: frame_vm_group_bin_12025 (RW)
0x1cf: frame_vm_group_bin_11901 (RW)
0x1d0: frame_vm_group_bin_21016 (RW)
0x1d1: frame_vm_group_bin_13843 (RW)
0x1d2: frame_vm_group_bin_6659 (RW)
0x1d3: frame_vm_group_bin_22855 (RW)
0x1d4: frame_vm_group_bin_15672 (RW)
0x1d5: frame_vm_group_bin_8482 (RW)
0x1d6: frame_vm_group_bin_1290 (RW)
0x1d7: frame_vm_group_bin_17480 (RW)
0x1d8: frame_vm_group_bin_10315 (RW)
0x1d9: frame_vm_group_bin_3155 (RW)
0x1d: frame_vm_group_bin_16393 (RW)
0x1da: frame_vm_group_bin_19225 (RW)
0x1db: frame_vm_group_bin_12054 (RW)
0x1dc: frame_vm_group_bin_16625 (RW)
0x1dd: frame_vm_group_bin_21051 (RW)
0x1de: frame_vm_group_bin_13874 (RW)
0x1df: frame_vm_group_bin_6693 (RW)
0x1e0: frame_vm_group_bin_22889 (RW)
0x1e1: frame_vm_group_bin_15706 (RW)
0x1e2: frame_vm_group_bin_8515 (RW)
0x1e3: frame_vm_group_bin_1323 (RW)
0x1e4: frame_vm_group_bin_17503 (RW)
0x1e5: frame_vm_group_bin_10349 (RW)
0x1e6: frame_vm_group_bin_3189 (RW)
0x1e7: frame_vm_group_bin_19258 (RW)
0x1e8: frame_vm_group_bin_12085 (RW)
0x1e9: frame_vm_group_bin_4986 (RW)
0x1e: frame_vm_group_bin_9212 (RW)
0x1ea: frame_vm_group_bin_21084 (RW)
0x1eb: frame_vm_group_bin_13906 (RW)
0x1ec: frame_vm_group_bin_6725 (RW)
0x1ed: frame_vm_group_bin_22922 (RW)
0x1ee: frame_vm_group_bin_15739 (RW)
0x1ef: frame_vm_group_bin_8547 (RW)
0x1f0: frame_vm_group_bin_1356 (RW)
0x1f1: frame_vm_group_bin_17531 (RW)
0x1f2: frame_vm_group_bin_10381 (RW)
0x1f3: frame_vm_group_bin_3222 (RW)
0x1f4: frame_vm_group_bin_19291 (RW)
0x1f5: frame_vm_group_bin_12117 (RW)
0x1f6: frame_vm_group_bin_5019 (RW)
0x1f7: frame_vm_group_bin_21117 (RW)
0x1f8: frame_vm_group_bin_13939 (RW)
0x1f9: frame_vm_group_bin_6757 (RW)
0x1f: frame_vm_group_bin_2030 (RW)
0x1fa: frame_vm_group_bin_22955 (RW)
0x1fb: frame_vm_group_bin_15773 (RW)
0x1fc: frame_vm_group_bin_8580 (RW)
0x1fd: frame_vm_group_bin_1391 (RW)
0x1fe: frame_vm_group_bin_14457 (RW)
0x1ff: frame_vm_group_bin_10409 (RW)
0x20: frame_vm_group_bin_18126 (RW)
0x21: frame_vm_group_bin_11038 (RW)
0x22: frame_vm_group_bin_3853 (RW)
0x23: frame_vm_group_bin_19951 (RW)
0x24: frame_vm_group_bin_12750 (RW)
0x25: frame_vm_group_bin_5686 (RW)
0x26: frame_vm_group_bin_21785 (RW)
0x27: frame_vm_group_bin_14611 (RW)
0x28: frame_vm_group_bin_7397 (RW)
0x29: frame_vm_group_bin_0256 (RW)
0x2: frame_vm_group_bin_0172 (RW)
0x2a: frame_vm_group_bin_16426 (RW)
0x2b: frame_vm_group_bin_9236 (RW)
0x2c: frame_vm_group_bin_2063 (RW)
0x2d: frame_vm_group_bin_18159 (RW)
0x2e: frame_vm_group_bin_11071 (RW)
0x2f: frame_vm_group_bin_3886 (RW)
0x30: frame_vm_group_bin_19984 (RW)
0x31: frame_vm_group_bin_12783 (RW)
0x32: frame_vm_group_bin_5719 (RW)
0x33: frame_vm_group_bin_21819 (RW)
0x34: frame_vm_group_bin_14644 (RW)
0x35: frame_vm_group_bin_7430 (RW)
0x36: frame_vm_group_bin_0280 (RW)
0x37: frame_vm_group_bin_16459 (RW)
0x38: frame_vm_group_bin_9259 (RW)
0x39: frame_vm_group_bin_2096 (RW)
0x3: frame_vm_group_bin_16326 (RW)
0x3a: frame_vm_group_bin_18192 (RW)
0x3b: frame_vm_group_bin_11105 (RW)
0x3c: frame_vm_group_bin_3920 (RW)
0x3d: frame_vm_group_bin_20016 (RW)
0x3e: frame_vm_group_bin_4292 (RW)
0x3f: frame_vm_group_bin_5749 (RW)
0x40: frame_vm_group_bin_21853 (RW)
0x41: frame_vm_group_bin_14678 (RW)
0x42: frame_vm_group_bin_7464 (RW)
0x43: frame_vm_group_bin_0311 (RW)
0x44: frame_vm_group_bin_16493 (RW)
0x45: frame_vm_group_bin_9285 (RW)
0x46: frame_vm_group_bin_2131 (RW)
0x47: frame_vm_group_bin_18225 (RW)
0x48: frame_vm_group_bin_11137 (RW)
0x49: frame_vm_group_bin_3952 (RW)
0x4: frame_vm_group_bin_9151 (RW)
0x4a: frame_vm_group_bin_20049 (RW)
0x4b: frame_vm_group_bin_12849 (RW)
0x4c: frame_vm_group_bin_5772 (RW)
0x4d: frame_vm_group_bin_21886 (RW)
0x4e: frame_vm_group_bin_14711 (RW)
0x4f: frame_vm_group_bin_7497 (RW)
0x50: frame_vm_group_bin_0343 (RW)
0x51: frame_vm_group_bin_16526 (RW)
0x52: frame_vm_group_bin_9314 (RW)
0x53: frame_vm_group_bin_2164 (RW)
0x54: frame_vm_group_bin_18258 (RW)
0x55: frame_vm_group_bin_11170 (RW)
0x56: frame_vm_group_bin_3985 (RW)
0x57: frame_vm_group_bin_20082 (RW)
0x58: frame_vm_group_bin_12882 (RW)
0x59: frame_vm_group_bin_5797 (RW)
0x5: frame_vm_group_bin_1963 (RW)
0x5a: frame_vm_group_bin_21919 (RW)
0x5b: frame_vm_group_bin_14744 (RW)
0x5c: frame_vm_group_bin_7831 (RW)
0x5d: frame_vm_group_bin_0375 (RW)
0x5e: frame_vm_group_bin_16559 (RW)
0x5f: frame_vm_group_bin_9348 (RW)
0x60: frame_vm_group_bin_2197 (RW)
0x61: frame_vm_group_bin_18292 (RW)
0x62: frame_vm_group_bin_11204 (RW)
0x63: frame_vm_group_bin_4019 (RW)
0x64: frame_vm_group_bin_20115 (RW)
0x65: frame_vm_group_bin_12916 (RW)
0x66: frame_vm_group_bin_5817 (RW)
0x67: frame_vm_group_bin_21952 (RW)
0x68: frame_vm_group_bin_13940 (RW)
0x69: frame_vm_group_bin_7561 (RW)
0x6: frame_vm_group_bin_18061 (RW)
0x6a: frame_vm_group_bin_0405 (RW)
0x6b: frame_vm_group_bin_16592 (RW)
0x6c: frame_vm_group_bin_9381 (RW)
0x6d: frame_vm_group_bin_2226 (RW)
0x6e: frame_vm_group_bin_18325 (RW)
0x6f: frame_vm_group_bin_11237 (RW)
0x70: frame_vm_group_bin_4052 (RW)
0x71: frame_vm_group_bin_20148 (RW)
0x72: frame_vm_group_bin_12948 (RW)
0x73: frame_vm_group_bin_5842 (RW)
0x74: frame_vm_group_bin_21985 (RW)
0x75: frame_vm_group_bin_14809 (RW)
0x76: frame_vm_group_bin_7594 (RW)
0x77: frame_vm_group_bin_0434 (RW)
0x78: frame_vm_group_bin_16624 (RW)
0x79: frame_vm_group_bin_9415 (RW)
0x7: frame_vm_group_bin_10971 (RW)
0x7a: frame_vm_group_bin_2256 (RW)
0x7b: frame_vm_group_bin_18359 (RW)
0x7c: frame_vm_group_bin_11271 (RW)
0x7d: frame_vm_group_bin_4086 (RW)
0x7e: frame_vm_group_bin_5761 (RW)
0x7f: frame_vm_group_bin_12982 (RW)
0x80: frame_vm_group_bin_5866 (RW)
0x81: frame_vm_group_bin_1387 (RW)
0x82: frame_vm_group_bin_14843 (RW)
0x83: frame_vm_group_bin_7628 (RW)
0x84: frame_vm_group_bin_0468 (RW)
0x85: frame_vm_group_bin_16658 (RW)
0x86: frame_vm_group_bin_9449 (RW)
0x87: frame_vm_group_bin_2289 (RW)
0x88: frame_vm_group_bin_14695 (RW)
0x89: frame_vm_group_bin_11304 (RW)
0x8: frame_vm_group_bin_3786 (RW)
0x8a: frame_vm_group_bin_4118 (RW)
0x8b: frame_vm_group_bin_20213 (RW)
0x8c: frame_vm_group_bin_13017 (RW)
0x8d: frame_vm_group_bin_5892 (RW)
0x8e: frame_vm_group_bin_6052 (RW)
0x8f: frame_vm_group_bin_14876 (RW)
0x90: frame_vm_group_bin_7661 (RW)
0x91: frame_vm_group_bin_0500 (RW)
0x92: frame_vm_group_bin_16691 (RW)
0x93: frame_vm_group_bin_9482 (RW)
0x94: frame_vm_group_bin_2322 (RW)
0x95: frame_vm_group_bin_18423 (RW)
0x96: frame_vm_group_bin_11337 (RW)
0x97: frame_vm_group_bin_4151 (RW)
0x98: frame_vm_group_bin_20246 (RW)
0x99: frame_vm_group_bin_13050 (RW)
0x9: frame_vm_group_bin_19886 (RW)
0x9a: frame_vm_group_bin_5919 (RW)
0x9b: frame_vm_group_bin_22065 (RW)
0x9c: frame_vm_group_bin_14910 (RW)
0x9d: frame_vm_group_bin_7695 (RW)
0x9e: frame_vm_group_bin_0533 (RW)
0x9f: frame_vm_group_bin_16725 (RW)
0xa0: frame_vm_group_bin_9516 (RW)
0xa1: frame_vm_group_bin_2356 (RW)
0xa2: frame_vm_group_bin_8672 (RW)
0xa3: frame_vm_group_bin_11369 (RW)
0xa4: frame_vm_group_bin_4184 (RW)
0xa5: frame_vm_group_bin_20279 (RW)
0xa6: frame_vm_group_bin_13084 (RW)
0xa7: frame_vm_group_bin_5942 (RW)
0xa8: frame_vm_group_bin_22093 (RW)
0xa9: frame_vm_group_bin_14943 (RW)
0xa: frame_vm_group_bin_12697 (RW)
0xaa: frame_vm_group_bin_7727 (RW)
0xab: frame_vm_group_bin_0564 (RW)
0xac: frame_vm_group_bin_16758 (RW)
0xad: frame_vm_group_bin_9549 (RW)
0xae: frame_vm_group_bin_2389 (RW)
0xaf: frame_vm_group_bin_5421 (RW)
0xb0: frame_vm_group_bin_11401 (RW)
0xb1: frame_vm_group_bin_4216 (RW)
0xb2: frame_vm_group_bin_20312 (RW)
0xb3: frame_vm_group_bin_13117 (RW)
0xb4: frame_vm_group_bin_5967 (RW)
0xb5: frame_vm_group_bin_22125 (RW)
0xb6: frame_vm_group_bin_14976 (RW)
0xb7: frame_vm_group_bin_7760 (RW)
0xb8: frame_vm_group_bin_0596 (RW)
0xb9: frame_vm_group_bin_16791 (RW)
0xb: frame_vm_group_bin_5619 (RW)
0xba: frame_vm_group_bin_9583 (RW)
0xbb: frame_vm_group_bin_11526 (RW)
0xbc: frame_vm_group_bin_18513 (RW)
0xbd: frame_vm_group_bin_11434 (RW)
0xbe: frame_vm_group_bin_4250 (RW)
0xbf: frame_vm_group_bin_20348 (RW)
0xc0: frame_vm_group_bin_13151 (RW)
0xc1: frame_vm_group_bin_5996 (RW)
0xc2: frame_vm_group_bin_22159 (RW)
0xc3: frame_vm_group_bin_15010 (RW)
0xc4: frame_vm_group_bin_7794 (RW)
0xc5: frame_vm_group_bin_0628 (RW)
0xc6: frame_vm_group_bin_16825 (RW)
0xc7: frame_vm_group_bin_9616 (RW)
0xc8: frame_vm_group_bin_2455 (RW)
0xc9: frame_vm_group_bin_18538 (RW)
0xc: frame_vm_group_bin_21719 (RW)
0xca: frame_vm_group_bin_11467 (RW)
0xcb: frame_vm_group_bin_4283 (RW)
0xcc: frame_vm_group_bin_20381 (RW)
0xcd: frame_vm_group_bin_13184 (RW)
0xce: frame_vm_group_bin_6027 (RW)
0xcf: frame_vm_group_bin_22192 (RW)
0xd0: frame_vm_group_bin_4694 (RW)
0xd1: frame_vm_group_bin_7827 (RW)
0xd2: frame_vm_group_bin_0662 (RW)
0xd3: frame_vm_group_bin_16858 (RW)
0xd4: frame_vm_group_bin_9649 (RW)
0xd5: frame_vm_group_bin_2487 (RW)
0xd6: frame_vm_group_bin_18564 (RW)
0xd7: frame_vm_group_bin_11500 (RW)
0xd8: frame_vm_group_bin_4316 (RW)
0xd9: frame_vm_group_bin_20414 (RW)
0xd: frame_vm_group_bin_14545 (RW)
0xda: frame_vm_group_bin_13218 (RW)
0xdb: frame_vm_group_bin_6054 (RW)
0xdc: frame_vm_group_bin_22226 (RW)
0xdd: frame_vm_group_bin_15066 (RW)
0xde: frame_vm_group_bin_7860 (RW)
0xdf: frame_vm_group_bin_0696 (RW)
0xe0: frame_vm_group_bin_16890 (RW)
0xe1: frame_vm_group_bin_9682 (RW)
0xe2: frame_vm_group_bin_2521 (RW)
0xe3: frame_vm_group_bin_18598 (RW)
0xe4: frame_vm_group_bin_11534 (RW)
0xe5: frame_vm_group_bin_4352 (RW)
0xe6: frame_vm_group_bin_20448 (RW)
0xe7: frame_vm_group_bin_13251 (RW)
0xe8: frame_vm_group_bin_6079 (RW)
0xe9: frame_vm_group_bin_22259 (RW)
0xe: frame_vm_group_bin_7330 (RW)
0xea: frame_vm_group_bin_15090 (RW)
0xeb: frame_vm_group_bin_7893 (RW)
0xec: frame_vm_group_bin_0729 (RW)
0xed: frame_vm_group_bin_16923 (RW)
0xee: frame_vm_group_bin_9715 (RW)
0xef: frame_vm_group_bin_2554 (RW)
0xf0: frame_vm_group_bin_18631 (RW)
0xf1: frame_vm_group_bin_11564 (RW)
0xf2: frame_vm_group_bin_4385 (RW)
0xf3: frame_vm_group_bin_20481 (RW)
0xf4: frame_vm_group_bin_13284 (RW)
0xf5: frame_vm_group_bin_6110 (RW)
0xf6: frame_vm_group_bin_22291 (RW)
0xf7: frame_vm_group_bin_15117 (RW)
0xf8: frame_vm_group_bin_7926 (RW)
0xf9: frame_vm_group_bin_0762 (RW)
0xf: frame_vm_group_bin_0204 (RW)
0xfa: frame_vm_group_bin_16957 (RW)
0xfb: frame_vm_group_bin_9749 (RW)
0xfc: frame_vm_group_bin_2588 (RW)
0xfd: frame_vm_group_bin_18664 (RW)
0xfe: frame_vm_group_bin_11593 (RW)
0xff: frame_vm_group_bin_4419 (RW)
}
pt_vm_group_bin_0220 {
0x0: frame_vm_group_bin_12656 (RW)
0x100: frame_vm_group_bin_18640 (RW)
0x101: frame_vm_group_bin_11574 (RW)
0x102: frame_vm_group_bin_4395 (RW)
0x103: frame_vm_group_bin_20491 (RW)
0x104: frame_vm_group_bin_13294 (RW)
0x105: frame_vm_group_bin_6119 (RW)
0x106: frame_vm_group_bin_22301 (RW)
0x107: frame_vm_group_bin_15126 (RW)
0x108: frame_vm_group_bin_7937 (RW)
0x109: frame_vm_group_bin_0772 (RW)
0x10: frame_vm_group_bin_14521 (RW)
0x10a: frame_vm_group_bin_16966 (RW)
0x10b: frame_vm_group_bin_9758 (RW)
0x10c: frame_vm_group_bin_2597 (RW)
0x10d: frame_vm_group_bin_18673 (RW)
0x10e: frame_vm_group_bin_11599 (RW)
0x10f: frame_vm_group_bin_4428 (RW)
0x110: frame_vm_group_bin_20524 (RW)
0x111: frame_vm_group_bin_13326 (RW)
0x112: frame_vm_group_bin_6151 (RW)
0x113: frame_vm_group_bin_22334 (RW)
0x114: frame_vm_group_bin_15149 (RW)
0x115: frame_vm_group_bin_7970 (RW)
0x116: frame_vm_group_bin_0805 (RW)
0x117: frame_vm_group_bin_16999 (RW)
0x118: frame_vm_group_bin_9791 (RW)
0x119: frame_vm_group_bin_2630 (RW)
0x11: frame_vm_group_bin_7306 (RW)
0x11a: frame_vm_group_bin_18706 (RW)
0x11b: frame_vm_group_bin_11627 (RW)
0x11c: frame_vm_group_bin_4462 (RW)
0x11d: frame_vm_group_bin_20558 (RW)
0x11e: frame_vm_group_bin_13360 (RW)
0x11f: frame_vm_group_bin_19552 (RW)
0x120: frame_vm_group_bin_22367 (RW)
0x121: frame_vm_group_bin_15183 (RW)
0x122: frame_vm_group_bin_8002 (RW)
0x123: frame_vm_group_bin_0838 (RW)
0x124: frame_vm_group_bin_17033 (RW)
0x125: frame_vm_group_bin_9825 (RW)
0x126: frame_vm_group_bin_2664 (RW)
0x127: frame_vm_group_bin_18737 (RW)
0x128: frame_vm_group_bin_11648 (RW)
0x129: frame_vm_group_bin_4495 (RW)
0x12: frame_vm_group_bin_0181 (RW)
0x12a: frame_vm_group_bin_20591 (RW)
0x12b: frame_vm_group_bin_13391 (RW)
0x12c: frame_vm_group_bin_0928 (RW)
0x12d: frame_vm_group_bin_22400 (RW)
0x12e: frame_vm_group_bin_15216 (RW)
0x12f: frame_vm_group_bin_8030 (RW)
0x130: frame_vm_group_bin_0871 (RW)
0x131: frame_vm_group_bin_17066 (RW)
0x132: frame_vm_group_bin_9858 (RW)
0x133: frame_vm_group_bin_2697 (RW)
0x134: frame_vm_group_bin_18770 (RW)
0x135: frame_vm_group_bin_11384 (RW)
0x136: frame_vm_group_bin_4528 (RW)
0x137: frame_vm_group_bin_20624 (RW)
0x138: frame_vm_group_bin_13424 (RW)
0x139: frame_vm_group_bin_6241 (RW)
0x13: frame_vm_group_bin_16335 (RW)
0x13a: frame_vm_group_bin_22433 (RW)
0x13b: frame_vm_group_bin_15251 (RW)
0x13c: frame_vm_group_bin_8061 (RW)
0x13d: frame_vm_group_bin_0905 (RW)
0x13e: frame_vm_group_bin_17100 (RW)
0x13f: frame_vm_group_bin_9891 (RW)
0x140: frame_vm_group_bin_2731 (RW)
0x141: frame_vm_group_bin_18804 (RW)
0x142: frame_vm_group_bin_16032 (RW)
0x143: frame_vm_group_bin_4561 (RW)
0x144: frame_vm_group_bin_20657 (RW)
0x145: frame_vm_group_bin_13458 (RW)
0x146: frame_vm_group_bin_6273 (RW)
0x147: frame_vm_group_bin_22466 (RW)
0x148: frame_vm_group_bin_15283 (RW)
0x149: frame_vm_group_bin_8093 (RW)
0x14: frame_vm_group_bin_9160 (RW)
0x14a: frame_vm_group_bin_0938 (RW)
0x14b: frame_vm_group_bin_17133 (RW)
0x14c: frame_vm_group_bin_9924 (RW)
0x14d: frame_vm_group_bin_2764 (RW)
0x14e: frame_vm_group_bin_18838 (RW)
0x14f: frame_vm_group_bin_20673 (RW)
0x150: frame_vm_group_bin_4586 (RW)
0x151: frame_vm_group_bin_20690 (RW)
0x152: frame_vm_group_bin_13491 (RW)
0x153: frame_vm_group_bin_6306 (RW)
0x154: frame_vm_group_bin_22499 (RW)
0x155: frame_vm_group_bin_15316 (RW)
0x156: frame_vm_group_bin_8125 (RW)
0x157: frame_vm_group_bin_0971 (RW)
0x158: frame_vm_group_bin_17165 (RW)
0x159: frame_vm_group_bin_9955 (RW)
0x15: frame_vm_group_bin_1972 (RW)
0x15a: frame_vm_group_bin_2798 (RW)
0x15b: frame_vm_group_bin_18872 (RW)
0x15c: frame_vm_group_bin_2024 (RW)
0x15d: frame_vm_group_bin_4610 (RW)
0x15e: frame_vm_group_bin_20724 (RW)
0x15f: frame_vm_group_bin_13525 (RW)
0x160: frame_vm_group_bin_6339 (RW)
0x161: frame_vm_group_bin_22532 (RW)
0x162: frame_vm_group_bin_15350 (RW)
0x163: frame_vm_group_bin_8159 (RW)
0x164: frame_vm_group_bin_1005 (RW)
0x165: frame_vm_group_bin_17196 (RW)
0x166: frame_vm_group_bin_9989 (RW)
0x167: frame_vm_group_bin_2831 (RW)
0x168: frame_vm_group_bin_18905 (RW)
0x169: frame_vm_group_bin_6663 (RW)
0x16: frame_vm_group_bin_18070 (RW)
0x16a: frame_vm_group_bin_4636 (RW)
0x16b: frame_vm_group_bin_20757 (RW)
0x16c: frame_vm_group_bin_13558 (RW)
0x16d: frame_vm_group_bin_0951 (RW)
0x16e: frame_vm_group_bin_22565 (RW)
0x16f: frame_vm_group_bin_15383 (RW)
0x170: frame_vm_group_bin_8192 (RW)
0x171: frame_vm_group_bin_1030 (RW)
0x172: frame_vm_group_bin_17229 (RW)
0x173: frame_vm_group_bin_10022 (RW)
0x174: frame_vm_group_bin_2863 (RW)
0x175: frame_vm_group_bin_18938 (RW)
0x176: frame_vm_group_bin_11795 (RW)
0x177: frame_vm_group_bin_4669 (RW)
0x178: frame_vm_group_bin_20790 (RW)
0x179: frame_vm_group_bin_13591 (RW)
0x17: frame_vm_group_bin_10980 (RW)
0x17a: frame_vm_group_bin_6403 (RW)
0x17b: frame_vm_group_bin_22599 (RW)
0x17c: frame_vm_group_bin_15417 (RW)
0x17d: frame_vm_group_bin_8226 (RW)
0x17e: frame_vm_group_bin_1053 (RW)
0x17f: frame_vm_group_bin_17262 (RW)
0x180: frame_vm_group_bin_10056 (RW)
0x181: frame_vm_group_bin_2899 (RW)
0x182: frame_vm_group_bin_17481 (RW)
0x183: frame_vm_group_bin_11828 (RW)
0x184: frame_vm_group_bin_4701 (RW)
0x185: frame_vm_group_bin_20823 (RW)
0x186: frame_vm_group_bin_13625 (RW)
0x187: frame_vm_group_bin_6435 (RW)
0x188: frame_vm_group_bin_22632 (RW)
0x189: frame_vm_group_bin_15450 (RW)
0x18: frame_vm_group_bin_3795 (RW)
0x18a: frame_vm_group_bin_8259 (RW)
0x18b: frame_vm_group_bin_1076 (RW)
0x18c: frame_vm_group_bin_17295 (RW)
0x18d: frame_vm_group_bin_10089 (RW)
0x18e: frame_vm_group_bin_2932 (RW)
0x18f: frame_vm_group_bin_19002 (RW)
0x190: frame_vm_group_bin_20698 (RW)
0x191: frame_vm_group_bin_4733 (RW)
0x192: frame_vm_group_bin_20852 (RW)
0x193: frame_vm_group_bin_13657 (RW)
0x194: frame_vm_group_bin_6468 (RW)
0x195: frame_vm_group_bin_22665 (RW)
0x196: frame_vm_group_bin_15483 (RW)
0x197: frame_vm_group_bin_8291 (RW)
0x198: frame_vm_group_bin_1103 (RW)
0x199: frame_vm_group_bin_17328 (RW)
0x19: frame_vm_group_bin_19895 (RW)
0x19a: frame_vm_group_bin_10123 (RW)
0x19b: frame_vm_group_bin_2966 (RW)
0x19c: frame_vm_group_bin_19036 (RW)
0x19d: frame_vm_group_bin_11887 (RW)
0x19e: frame_vm_group_bin_4767 (RW)
0x19f: frame_vm_group_bin_20878 (RW)
0x1: frame_vm_group_bin_5565 (RW)
0x1a0: frame_vm_group_bin_13691 (RW)
0x1a1: frame_vm_group_bin_6502 (RW)
0x1a2: frame_vm_group_bin_22699 (RW)
0x1a3: frame_vm_group_bin_15516 (RW)
0x1a4: frame_vm_group_bin_8325 (RW)
0x1a5: frame_vm_group_bin_1136 (RW)
0x1a6: frame_vm_group_bin_17361 (RW)
0x1a7: frame_vm_group_bin_10158 (RW)
0x1a8: frame_vm_group_bin_2999 (RW)
0x1a9: frame_vm_group_bin_19069 (RW)
0x1a: frame_vm_group_bin_12705 (RW)
0x1aa: frame_vm_group_bin_11910 (RW)
0x1ab: frame_vm_group_bin_4800 (RW)
0x1ac: frame_vm_group_bin_20905 (RW)
0x1ad: frame_vm_group_bin_13723 (RW)
0x1ae: frame_vm_group_bin_6535 (RW)
0x1af: frame_vm_group_bin_22732 (RW)
0x1b0: frame_vm_group_bin_15548 (RW)
0x1b1: frame_vm_group_bin_8358 (RW)
0x1b2: frame_vm_group_bin_1169 (RW)
0x1b3: frame_vm_group_bin_17391 (RW)
0x1b4: frame_vm_group_bin_10191 (RW)
0x1b5: frame_vm_group_bin_3032 (RW)
0x1b6: frame_vm_group_bin_19102 (RW)
0x1b7: frame_vm_group_bin_11430 (RW)
0x1b8: frame_vm_group_bin_4832 (RW)
0x1b9: frame_vm_group_bin_20933 (RW)
0x1b: frame_vm_group_bin_5629 (RW)
0x1ba: frame_vm_group_bin_13758 (RW)
0x1bb: frame_vm_group_bin_6569 (RW)
0x1bc: frame_vm_group_bin_22765 (RW)
0x1bd: frame_vm_group_bin_15582 (RW)
0x1be: frame_vm_group_bin_8392 (RW)
0x1bf: frame_vm_group_bin_1203 (RW)
0x1c0: frame_vm_group_bin_17419 (RW)
0x1c1: frame_vm_group_bin_10225 (RW)
0x1c2: frame_vm_group_bin_3066 (RW)
0x1c3: frame_vm_group_bin_19134 (RW)
0x1c4: frame_vm_group_bin_11971 (RW)
0x1c5: frame_vm_group_bin_4866 (RW)
0x1c6: frame_vm_group_bin_20961 (RW)
0x1c7: frame_vm_group_bin_13791 (RW)
0x1c8: frame_vm_group_bin_6602 (RW)
0x1c9: frame_vm_group_bin_22798 (RW)
0x1c: frame_vm_group_bin_21729 (RW)
0x1ca: frame_vm_group_bin_15615 (RW)
0x1cb: frame_vm_group_bin_8425 (RW)
0x1cc: frame_vm_group_bin_1236 (RW)
0x1cd: frame_vm_group_bin_17444 (RW)
0x1ce: frame_vm_group_bin_10258 (RW)
0x1cf: frame_vm_group_bin_3099 (RW)
0x1d0: frame_vm_group_bin_19167 (RW)
0x1d1: frame_vm_group_bin_12003 (RW)
0x1d2: frame_vm_group_bin_4899 (RW)
0x1d3: frame_vm_group_bin_20992 (RW)
0x1d4: frame_vm_group_bin_13822 (RW)
0x1d5: frame_vm_group_bin_6635 (RW)
0x1d6: frame_vm_group_bin_22831 (RW)
0x1d7: frame_vm_group_bin_15648 (RW)
0x1d8: frame_vm_group_bin_8458 (RW)
0x1d9: frame_vm_group_bin_1268 (RW)
0x1d: frame_vm_group_bin_14555 (RW)
0x1da: frame_vm_group_bin_7786 (RW)
0x1db: frame_vm_group_bin_10292 (RW)
0x1dc: frame_vm_group_bin_3132 (RW)
0x1dd: frame_vm_group_bin_19201 (RW)
0x1de: frame_vm_group_bin_12034 (RW)
0x1df: frame_vm_group_bin_4931 (RW)
0x1e0: frame_vm_group_bin_21026 (RW)
0x1e1: frame_vm_group_bin_13853 (RW)
0x1e2: frame_vm_group_bin_6669 (RW)
0x1e3: frame_vm_group_bin_22865 (RW)
0x1e4: frame_vm_group_bin_15682 (RW)
0x1e5: frame_vm_group_bin_8492 (RW)
0x1e6: frame_vm_group_bin_1300 (RW)
0x1e7: frame_vm_group_bin_17487 (RW)
0x1e8: frame_vm_group_bin_10325 (RW)
0x1e9: frame_vm_group_bin_3165 (RW)
0x1e: frame_vm_group_bin_7340 (RW)
0x1ea: frame_vm_group_bin_19234 (RW)
0x1eb: frame_vm_group_bin_6710 (RW)
0x1ec: frame_vm_group_bin_4963 (RW)
0x1ed: frame_vm_group_bin_21060 (RW)
0x1ee: frame_vm_group_bin_13882 (RW)
0x1ef: frame_vm_group_bin_6702 (RW)
0x1f0: frame_vm_group_bin_22898 (RW)
0x1f1: frame_vm_group_bin_15715 (RW)
0x1f2: frame_vm_group_bin_8524 (RW)
0x1f3: frame_vm_group_bin_1332 (RW)
0x1f4: frame_vm_group_bin_17511 (RW)
0x1f5: frame_vm_group_bin_10358 (RW)
0x1f6: frame_vm_group_bin_3198 (RW)
0x1f7: frame_vm_group_bin_19267 (RW)
0x1f8: frame_vm_group_bin_12094 (RW)
0x1f9: frame_vm_group_bin_4995 (RW)
0x1f: frame_vm_group_bin_13733 (RW)
0x1fa: frame_vm_group_bin_21094 (RW)
0x1fb: frame_vm_group_bin_13916 (RW)
0x1fc: frame_vm_group_bin_6735 (RW)
0x1fd: frame_vm_group_bin_22932 (RW)
0x1fe: frame_vm_group_bin_15749 (RW)
0x1ff: frame_vm_group_bin_8556 (RW)
0x20: frame_vm_group_bin_16369 (RW)
0x21: frame_vm_group_bin_9192 (RW)
0x22: frame_vm_group_bin_2006 (RW)
0x23: frame_vm_group_bin_18102 (RW)
0x24: frame_vm_group_bin_11014 (RW)
0x25: frame_vm_group_bin_3829 (RW)
0x26: frame_vm_group_bin_19927 (RW)
0x27: frame_vm_group_bin_12731 (RW)
0x28: frame_vm_group_bin_5662 (RW)
0x29: frame_vm_group_bin_21762 (RW)
0x2: frame_vm_group_bin_21663 (RW)
0x2a: frame_vm_group_bin_14588 (RW)
0x2b: frame_vm_group_bin_7373 (RW)
0x2c: frame_vm_group_bin_18380 (RW)
0x2d: frame_vm_group_bin_16402 (RW)
0x2e: frame_vm_group_bin_9219 (RW)
0x2f: frame_vm_group_bin_2039 (RW)
0x30: frame_vm_group_bin_18135 (RW)
0x31: frame_vm_group_bin_11047 (RW)
0x32: frame_vm_group_bin_3862 (RW)
0x33: frame_vm_group_bin_19960 (RW)
0x34: frame_vm_group_bin_12759 (RW)
0x35: frame_vm_group_bin_5695 (RW)
0x36: frame_vm_group_bin_21794 (RW)
0x37: frame_vm_group_bin_14620 (RW)
0x38: frame_vm_group_bin_7406 (RW)
0x39: frame_vm_group_bin_23119 (RW)
0x3: frame_vm_group_bin_14487 (RW)
0x3a: frame_vm_group_bin_16436 (RW)
0x3b: frame_vm_group_bin_9244 (RW)
0x3c: frame_vm_group_bin_2073 (RW)
0x3d: frame_vm_group_bin_18169 (RW)
0x3e: frame_vm_group_bin_11081 (RW)
0x3f: frame_vm_group_bin_3896 (RW)
0x40: frame_vm_group_bin_19992 (RW)
0x41: frame_vm_group_bin_12793 (RW)
0x42: frame_vm_group_bin_5729 (RW)
0x43: frame_vm_group_bin_21829 (RW)
0x44: frame_vm_group_bin_14654 (RW)
0x45: frame_vm_group_bin_7440 (RW)
0x46: frame_vm_group_bin_0289 (RW)
0x47: frame_vm_group_bin_16469 (RW)
0x48: frame_vm_group_bin_9267 (RW)
0x49: frame_vm_group_bin_2106 (RW)
0x4: frame_vm_group_bin_7274 (RW)
0x4a: frame_vm_group_bin_18201 (RW)
0x4b: frame_vm_group_bin_11114 (RW)
0x4c: frame_vm_group_bin_3929 (RW)
0x4d: frame_vm_group_bin_20025 (RW)
0x4e: frame_vm_group_bin_12825 (RW)
0x4f: frame_vm_group_bin_5755 (RW)
0x50: frame_vm_group_bin_21862 (RW)
0x51: frame_vm_group_bin_14687 (RW)
0x52: frame_vm_group_bin_7473 (RW)
0x53: frame_vm_group_bin_0320 (RW)
0x54: frame_vm_group_bin_16502 (RW)
0x55: frame_vm_group_bin_9293 (RW)
0x56: frame_vm_group_bin_2140 (RW)
0x57: frame_vm_group_bin_18234 (RW)
0x58: frame_vm_group_bin_11146 (RW)
0x59: frame_vm_group_bin_3961 (RW)
0x5: frame_vm_group_bin_4461 (RW)
0x5a: frame_vm_group_bin_20059 (RW)
0x5b: frame_vm_group_bin_12859 (RW)
0x5c: frame_vm_group_bin_5780 (RW)
0x5d: frame_vm_group_bin_21896 (RW)
0x5e: frame_vm_group_bin_14721 (RW)
0x5f: frame_vm_group_bin_7506 (RW)
0x60: frame_vm_group_bin_0352 (RW)
0x61: frame_vm_group_bin_16536 (RW)
0x62: frame_vm_group_bin_9324 (RW)
0x63: frame_vm_group_bin_2174 (RW)
0x64: frame_vm_group_bin_18268 (RW)
0x65: frame_vm_group_bin_11180 (RW)
0x66: frame_vm_group_bin_3995 (RW)
0x67: frame_vm_group_bin_20092 (RW)
0x68: frame_vm_group_bin_12892 (RW)
0x69: frame_vm_group_bin_5802 (RW)
0x6: frame_vm_group_bin_16303 (RW)
0x6a: frame_vm_group_bin_21928 (RW)
0x6b: frame_vm_group_bin_14753 (RW)
0x6c: frame_vm_group_bin_7538 (RW)
0x6d: frame_vm_group_bin_0384 (RW)
0x6e: frame_vm_group_bin_16568 (RW)
0x6f: frame_vm_group_bin_9357 (RW)
0x70: frame_vm_group_bin_2205 (RW)
0x71: frame_vm_group_bin_18301 (RW)
0x72: frame_vm_group_bin_11213 (RW)
0x73: frame_vm_group_bin_4028 (RW)
0x74: frame_vm_group_bin_20124 (RW)
0x75: frame_vm_group_bin_12925 (RW)
0x76: frame_vm_group_bin_5823 (RW)
0x77: frame_vm_group_bin_21961 (RW)
0x78: frame_vm_group_bin_14785 (RW)
0x79: frame_vm_group_bin_7570 (RW)
0x7: frame_vm_group_bin_9128 (RW)
0x7a: frame_vm_group_bin_0413 (RW)
0x7b: frame_vm_group_bin_16601 (RW)
0x7c: frame_vm_group_bin_9392 (RW)
0x7d: frame_vm_group_bin_2234 (RW)
0x7e: frame_vm_group_bin_18335 (RW)
0x7f: frame_vm_group_bin_11247 (RW)
0x80: frame_vm_group_bin_4062 (RW)
0x81: frame_vm_group_bin_20157 (RW)
0x82: frame_vm_group_bin_12958 (RW)
0x83: frame_vm_group_bin_10220 (RW)
0x84: frame_vm_group_bin_21995 (RW)
0x85: frame_vm_group_bin_14819 (RW)
0x86: frame_vm_group_bin_7604 (RW)
0x87: frame_vm_group_bin_0444 (RW)
0x88: frame_vm_group_bin_16634 (RW)
0x89: frame_vm_group_bin_9425 (RW)
0x8: frame_vm_group_bin_1940 (RW)
0x8a: frame_vm_group_bin_2265 (RW)
0x8b: frame_vm_group_bin_18368 (RW)
0x8c: frame_vm_group_bin_11280 (RW)
0x8d: frame_vm_group_bin_4095 (RW)
0x8e: frame_vm_group_bin_20189 (RW)
0x8f: frame_vm_group_bin_12991 (RW)
0x90: frame_vm_group_bin_5874 (RW)
0x91: frame_vm_group_bin_22024 (RW)
0x92: frame_vm_group_bin_14852 (RW)
0x93: frame_vm_group_bin_7637 (RW)
0x94: frame_vm_group_bin_0477 (RW)
0x95: frame_vm_group_bin_16667 (RW)
0x96: frame_vm_group_bin_9458 (RW)
0x97: frame_vm_group_bin_2298 (RW)
0x98: frame_vm_group_bin_18400 (RW)
0x99: frame_vm_group_bin_11313 (RW)
0x9: frame_vm_group_bin_18038 (RW)
0x9a: frame_vm_group_bin_4128 (RW)
0x9b: frame_vm_group_bin_20223 (RW)
0x9c: frame_vm_group_bin_13027 (RW)
0x9d: frame_vm_group_bin_5900 (RW)
0x9e: frame_vm_group_bin_22047 (RW)
0x9f: frame_vm_group_bin_14886 (RW)
0xa0: frame_vm_group_bin_7671 (RW)
0xa1: frame_vm_group_bin_0510 (RW)
0xa2: frame_vm_group_bin_16700 (RW)
0xa3: frame_vm_group_bin_9492 (RW)
0xa4: frame_vm_group_bin_2332 (RW)
0xa5: frame_vm_group_bin_18433 (RW)
0xa6: frame_vm_group_bin_11345 (RW)
0xa7: frame_vm_group_bin_4160 (RW)
0xa8: frame_vm_group_bin_20256 (RW)
0xa9: frame_vm_group_bin_13060 (RW)
0xa: frame_vm_group_bin_10948 (RW)
0xaa: frame_vm_group_bin_5927 (RW)
0xab: frame_vm_group_bin_22071 (RW)
0xac: frame_vm_group_bin_14919 (RW)
0xad: frame_vm_group_bin_7704 (RW)
0xae: frame_vm_group_bin_0542 (RW)
0xaf: frame_vm_group_bin_16734 (RW)
0xb0: frame_vm_group_bin_9525 (RW)
0xb1: frame_vm_group_bin_2365 (RW)
0xb2: frame_vm_group_bin_18464 (RW)
0xb3: frame_vm_group_bin_11378 (RW)
0xb4: frame_vm_group_bin_4193 (RW)
0xb5: frame_vm_group_bin_20288 (RW)
0xb6: frame_vm_group_bin_13093 (RW)
0xb7: frame_vm_group_bin_5606 (RW)
0xb8: frame_vm_group_bin_22101 (RW)
0xb9: frame_vm_group_bin_14952 (RW)
0xb: frame_vm_group_bin_3763 (RW)
0xba: frame_vm_group_bin_7737 (RW)
0xbb: frame_vm_group_bin_0574 (RW)
0xbc: frame_vm_group_bin_16768 (RW)
0xbd: frame_vm_group_bin_9559 (RW)
0xbe: frame_vm_group_bin_2399 (RW)
0xbf: frame_vm_group_bin_18493 (RW)
0xc0: frame_vm_group_bin_11410 (RW)
0xc1: frame_vm_group_bin_4226 (RW)
0xc2: frame_vm_group_bin_20324 (RW)
0xc3: frame_vm_group_bin_13127 (RW)
0xc4: frame_vm_group_bin_5974 (RW)
0xc5: frame_vm_group_bin_22135 (RW)
0xc6: frame_vm_group_bin_14986 (RW)
0xc7: frame_vm_group_bin_7770 (RW)
0xc8: frame_vm_group_bin_0606 (RW)
0xc9: frame_vm_group_bin_16801 (RW)
0xc: frame_vm_group_bin_19863 (RW)
0xca: frame_vm_group_bin_9592 (RW)
0xcb: frame_vm_group_bin_2431 (RW)
0xcc: frame_vm_group_bin_18520 (RW)
0xcd: frame_vm_group_bin_11443 (RW)
0xce: frame_vm_group_bin_4259 (RW)
0xcf: frame_vm_group_bin_20357 (RW)
0xd0: frame_vm_group_bin_13160 (RW)
0xd1: frame_vm_group_bin_6005 (RW)
0xd2: frame_vm_group_bin_22168 (RW)
0xd3: frame_vm_group_bin_15019 (RW)
0xd4: frame_vm_group_bin_7803 (RW)
0xd5: frame_vm_group_bin_0637 (RW)
0xd6: frame_vm_group_bin_16834 (RW)
0xd7: frame_vm_group_bin_9625 (RW)
0xd8: frame_vm_group_bin_2464 (RW)
0xd9: frame_vm_group_bin_18544 (RW)
0xd: frame_vm_group_bin_12680 (RW)
0xda: frame_vm_group_bin_11477 (RW)
0xdb: frame_vm_group_bin_4293 (RW)
0xdc: frame_vm_group_bin_20391 (RW)
0xdd: frame_vm_group_bin_13194 (RW)
0xde: frame_vm_group_bin_6037 (RW)
0xdf: frame_vm_group_bin_22202 (RW)
0xe0: frame_vm_group_bin_15048 (RW)
0xe1: frame_vm_group_bin_7836 (RW)
0xe2: frame_vm_group_bin_0672 (RW)
0xe3: frame_vm_group_bin_16867 (RW)
0xe4: frame_vm_group_bin_9659 (RW)
0xe5: frame_vm_group_bin_2497 (RW)
0xe6: frame_vm_group_bin_18574 (RW)
0xe7: frame_vm_group_bin_11510 (RW)
0xe8: frame_vm_group_bin_4326 (RW)
0xe9: frame_vm_group_bin_20424 (RW)
0xe: frame_vm_group_bin_5597 (RW)
0xea: frame_vm_group_bin_13227 (RW)
0xeb: frame_vm_group_bin_0904 (RW)
0xec: frame_vm_group_bin_22235 (RW)
0xed: frame_vm_group_bin_15072 (RW)
0xee: frame_vm_group_bin_7869 (RW)
0xef: frame_vm_group_bin_0705 (RW)
0xf0: frame_vm_group_bin_16899 (RW)
0xf1: frame_vm_group_bin_9691 (RW)
0xf2: frame_vm_group_bin_2530 (RW)
0xf3: frame_vm_group_bin_18607 (RW)
0xf4: frame_vm_group_bin_11543 (RW)
0xf5: frame_vm_group_bin_4361 (RW)
0xf6: frame_vm_group_bin_20457 (RW)
0xf7: frame_vm_group_bin_13260 (RW)
0xf8: frame_vm_group_bin_6088 (RW)
0xf9: frame_vm_group_bin_22268 (RW)
0xf: frame_vm_group_bin_21695 (RW)
0xfa: frame_vm_group_bin_15097 (RW)
0xfb: frame_vm_group_bin_7903 (RW)
0xfc: frame_vm_group_bin_0739 (RW)
0xfd: frame_vm_group_bin_16933 (RW)
0xfe: frame_vm_group_bin_9725 (RW)
0xff: frame_vm_group_bin_2564 (RW)
}
pt_vm_group_bin_0239 {
0x0: frame_vm_group_bin_15608 (RW)
0x100: frame_vm_group_bin_21615 (RW)
0x101: frame_vm_group_bin_14439 (RW)
0x102: frame_vm_group_bin_7226 (RW)
0x103: frame_vm_group_bin_13074 (RW)
0x104: frame_vm_group_bin_16260 (RW)
0x105: frame_vm_group_bin_9080 (RW)
0x106: frame_vm_group_bin_1892 (RW)
0x107: frame_vm_group_bin_17990 (RW)
0x108: frame_vm_group_bin_10900 (RW)
0x109: frame_vm_group_bin_3715 (RW)
0x10: frame_vm_group_bin_11920 (RW)
0x10a: frame_vm_group_bin_19815 (RW)
0x10b: frame_vm_group_bin_12642 (RW)
0x10c: frame_vm_group_bin_5550 (RW)
0x10d: frame_vm_group_bin_21648 (RW)
0x10e: frame_vm_group_bin_14472 (RW)
0x10f: frame_vm_group_bin_7259 (RW)
0x110: frame_vm_group_bin_17747 (RW)
0x111: frame_vm_group_bin_16289 (RW)
0x112: frame_vm_group_bin_9113 (RW)
0x113: frame_vm_group_bin_1925 (RW)
0x114: frame_vm_group_bin_18023 (RW)
0x115: frame_vm_group_bin_10933 (RW)
0x116: frame_vm_group_bin_3748 (RW)
0x117: frame_vm_group_bin_19848 (RW)
0x118: frame_vm_group_bin_12669 (RW)
0x119: frame_vm_group_bin_5582 (RW)
0x11: frame_vm_group_bin_10284 (RW)
0x11a: frame_vm_group_bin_21681 (RW)
0x11b: frame_vm_group_bin_14507 (RW)
0x11c: frame_vm_group_bin_7292 (RW)
0x11d: frame_vm_group_bin_22457 (RW)
0x11e: frame_vm_group_bin_16321 (RW)
0x11f: frame_vm_group_bin_9146 (RW)
0x120: frame_vm_group_bin_1958 (RW)
0x121: frame_vm_group_bin_18056 (RW)
0x122: frame_vm_group_bin_10966 (RW)
0x123: frame_vm_group_bin_3781 (RW)
0x124: frame_vm_group_bin_19881 (RW)
0x125: frame_vm_group_bin_12695 (RW)
0x126: frame_vm_group_bin_5614 (RW)
0x127: frame_vm_group_bin_21714 (RW)
0x128: frame_vm_group_bin_14540 (RW)
0x129: frame_vm_group_bin_7325 (RW)
0x12: frame_vm_group_bin_3124 (RW)
0x12a: frame_vm_group_bin_0199 (RW)
0x12b: frame_vm_group_bin_16354 (RW)
0x12c: frame_vm_group_bin_9178 (RW)
0x12d: frame_vm_group_bin_1991 (RW)
0x12e: frame_vm_group_bin_18088 (RW)
0x12f: frame_vm_group_bin_10999 (RW)
0x130: frame_vm_group_bin_3814 (RW)
0x131: frame_vm_group_bin_19913 (RW)
0x132: frame_vm_group_bin_12720 (RW)
0x133: frame_vm_group_bin_5647 (RW)
0x134: frame_vm_group_bin_21747 (RW)
0x135: frame_vm_group_bin_14573 (RW)
0x136: frame_vm_group_bin_7358 (RW)
0x137: frame_vm_group_bin_8460 (RW)
0x138: frame_vm_group_bin_16387 (RW)
0x139: frame_vm_group_bin_9206 (RW)
0x13: frame_vm_group_bin_19193 (RW)
0x13a: frame_vm_group_bin_2025 (RW)
0x13b: frame_vm_group_bin_18121 (RW)
0x13c: frame_vm_group_bin_11033 (RW)
0x13d: frame_vm_group_bin_3848 (RW)
0x13e: frame_vm_group_bin_19946 (RW)
0x13f: frame_vm_group_bin_12746 (RW)
0x140: frame_vm_group_bin_5681 (RW)
0x141: frame_vm_group_bin_21780 (RW)
0x142: frame_vm_group_bin_14606 (RW)
0x143: frame_vm_group_bin_7392 (RW)
0x144: frame_vm_group_bin_13097 (RW)
0x145: frame_vm_group_bin_16421 (RW)
0x146: frame_vm_group_bin_9234 (RW)
0x147: frame_vm_group_bin_2058 (RW)
0x148: frame_vm_group_bin_18154 (RW)
0x149: frame_vm_group_bin_11066 (RW)
0x14: frame_vm_group_bin_12027 (RW)
0x14a: frame_vm_group_bin_3881 (RW)
0x14b: frame_vm_group_bin_19979 (RW)
0x14c: frame_vm_group_bin_12778 (RW)
0x14d: frame_vm_group_bin_5714 (RW)
0x14e: frame_vm_group_bin_21814 (RW)
0x14f: frame_vm_group_bin_14639 (RW)
0x150: frame_vm_group_bin_7425 (RW)
0x151: frame_vm_group_bin_17768 (RW)
0x152: frame_vm_group_bin_16454 (RW)
0x153: frame_vm_group_bin_9257 (RW)
0x154: frame_vm_group_bin_2091 (RW)
0x155: frame_vm_group_bin_18187 (RW)
0x156: frame_vm_group_bin_11099 (RW)
0x157: frame_vm_group_bin_3914 (RW)
0x158: frame_vm_group_bin_20010 (RW)
0x159: frame_vm_group_bin_12811 (RW)
0x15: frame_vm_group_bin_4924 (RW)
0x15a: frame_vm_group_bin_5745 (RW)
0x15b: frame_vm_group_bin_21848 (RW)
0x15c: frame_vm_group_bin_14673 (RW)
0x15d: frame_vm_group_bin_7459 (RW)
0x15e: frame_vm_group_bin_0306 (RW)
0x15f: frame_vm_group_bin_16488 (RW)
0x160: frame_vm_group_bin_9283 (RW)
0x161: frame_vm_group_bin_2126 (RW)
0x162: frame_vm_group_bin_18220 (RW)
0x163: frame_vm_group_bin_11132 (RW)
0x164: frame_vm_group_bin_3947 (RW)
0x165: frame_vm_group_bin_20044 (RW)
0x166: frame_vm_group_bin_12844 (RW)
0x167: frame_vm_group_bin_5770 (RW)
0x168: frame_vm_group_bin_21881 (RW)
0x169: frame_vm_group_bin_14706 (RW)
0x16: frame_vm_group_bin_21018 (RW)
0x16a: frame_vm_group_bin_7492 (RW)
0x16b: frame_vm_group_bin_0338 (RW)
0x16c: frame_vm_group_bin_16521 (RW)
0x16d: frame_vm_group_bin_9310 (RW)
0x16e: frame_vm_group_bin_2159 (RW)
0x16f: frame_vm_group_bin_18253 (RW)
0x170: frame_vm_group_bin_11165 (RW)
0x171: frame_vm_group_bin_3980 (RW)
0x172: frame_vm_group_bin_20077 (RW)
0x173: frame_vm_group_bin_12877 (RW)
0x174: frame_vm_group_bin_5793 (RW)
0x175: frame_vm_group_bin_21914 (RW)
0x176: frame_vm_group_bin_14738 (RW)
0x177: frame_vm_group_bin_7524 (RW)
0x178: frame_vm_group_bin_8483 (RW)
0x179: frame_vm_group_bin_16553 (RW)
0x17: frame_vm_group_bin_13845 (RW)
0x17a: frame_vm_group_bin_9343 (RW)
0x17b: frame_vm_group_bin_2192 (RW)
0x17c: frame_vm_group_bin_18287 (RW)
0x17d: frame_vm_group_bin_11199 (RW)
0x17e: frame_vm_group_bin_4014 (RW)
0x17f: frame_vm_group_bin_20110 (RW)
0x180: frame_vm_group_bin_12911 (RW)
0x181: frame_vm_group_bin_18847 (RW)
0x182: frame_vm_group_bin_21947 (RW)
0x183: frame_vm_group_bin_14772 (RW)
0x184: frame_vm_group_bin_7556 (RW)
0x185: frame_vm_group_bin_13120 (RW)
0x186: frame_vm_group_bin_16587 (RW)
0x187: frame_vm_group_bin_9376 (RW)
0x188: frame_vm_group_bin_2222 (RW)
0x189: frame_vm_group_bin_18320 (RW)
0x18: frame_vm_group_bin_6661 (RW)
0x18a: frame_vm_group_bin_11232 (RW)
0x18b: frame_vm_group_bin_4047 (RW)
0x18c: frame_vm_group_bin_20143 (RW)
0x18d: frame_vm_group_bin_12943 (RW)
0x18e: frame_vm_group_bin_0246 (RW)
0x18f: frame_vm_group_bin_21980 (RW)
0x190: frame_vm_group_bin_14804 (RW)
0x191: frame_vm_group_bin_7589 (RW)
0x192: frame_vm_group_bin_0429 (RW)
0x193: frame_vm_group_bin_16619 (RW)
0x194: frame_vm_group_bin_9410 (RW)
0x195: frame_vm_group_bin_2250 (RW)
0x196: frame_vm_group_bin_18353 (RW)
0x197: frame_vm_group_bin_11265 (RW)
0x198: frame_vm_group_bin_4080 (RW)
0x199: frame_vm_group_bin_20175 (RW)
0x19: frame_vm_group_bin_22857 (RW)
0x19a: frame_vm_group_bin_12977 (RW)
0x19b: frame_vm_group_bin_4952 (RW)
0x19c: frame_vm_group_bin_22013 (RW)
0x19d: frame_vm_group_bin_14838 (RW)
0x19e: frame_vm_group_bin_7623 (RW)
0x19f: frame_vm_group_bin_0463 (RW)
0x1: frame_vm_group_bin_8418 (RW)
0x1a0: frame_vm_group_bin_16653 (RW)
0x1a1: frame_vm_group_bin_9444 (RW)
0x1a2: frame_vm_group_bin_2284 (RW)
0x1a3: frame_vm_group_bin_18387 (RW)
0x1a4: frame_vm_group_bin_11299 (RW)
0x1a5: frame_vm_group_bin_4113 (RW)
0x1a6: frame_vm_group_bin_20208 (RW)
0x1a7: frame_vm_group_bin_13012 (RW)
0x1a8: frame_vm_group_bin_5887 (RW)
0x1a9: frame_vm_group_bin_22039 (RW)
0x1a: frame_vm_group_bin_15675 (RW)
0x1aa: frame_vm_group_bin_14871 (RW)
0x1ab: frame_vm_group_bin_7656 (RW)
0x1ac: frame_vm_group_bin_0495 (RW)
0x1ad: frame_vm_group_bin_16686 (RW)
0x1ae: frame_vm_group_bin_9477 (RW)
0x1af: frame_vm_group_bin_2317 (RW)
0x1b0: frame_vm_group_bin_18418 (RW)
0x1b1: frame_vm_group_bin_11332 (RW)
0x1b2: frame_vm_group_bin_4146 (RW)
0x1b3: frame_vm_group_bin_20241 (RW)
0x1b4: frame_vm_group_bin_13045 (RW)
0x1b5: frame_vm_group_bin_14247 (RW)
0x1b6: frame_vm_group_bin_22060 (RW)
0x1b7: frame_vm_group_bin_14904 (RW)
0x1b8: frame_vm_group_bin_7689 (RW)
0x1b9: frame_vm_group_bin_0527 (RW)
0x1b: frame_vm_group_bin_8485 (RW)
0x1ba: frame_vm_group_bin_16720 (RW)
0x1bb: frame_vm_group_bin_9511 (RW)
0x1bc: frame_vm_group_bin_2351 (RW)
0x1bd: frame_vm_group_bin_18452 (RW)
0x1be: frame_vm_group_bin_11364 (RW)
0x1bf: frame_vm_group_bin_4179 (RW)
0x1c0: frame_vm_group_bin_20274 (RW)
0x1c1: frame_vm_group_bin_13079 (RW)
0x1c2: frame_vm_group_bin_18871 (RW)
0x1c3: frame_vm_group_bin_22089 (RW)
0x1c4: frame_vm_group_bin_14938 (RW)
0x1c5: frame_vm_group_bin_7722 (RW)
0x1c6: frame_vm_group_bin_0559 (RW)
0x1c7: frame_vm_group_bin_16753 (RW)
0x1c8: frame_vm_group_bin_9544 (RW)
0x1c9: frame_vm_group_bin_2384 (RW)
0x1c: frame_vm_group_bin_1293 (RW)
0x1ca: frame_vm_group_bin_18480 (RW)
0x1cb: frame_vm_group_bin_11396 (RW)
0x1cc: frame_vm_group_bin_4211 (RW)
0x1cd: frame_vm_group_bin_20307 (RW)
0x1ce: frame_vm_group_bin_13112 (RW)
0x1cf: frame_vm_group_bin_5962 (RW)
0x1d0: frame_vm_group_bin_22120 (RW)
0x1d1: frame_vm_group_bin_14971 (RW)
0x1d2: frame_vm_group_bin_7755 (RW)
0x1d3: frame_vm_group_bin_0591 (RW)
0x1d4: frame_vm_group_bin_16786 (RW)
0x1d5: frame_vm_group_bin_9577 (RW)
0x1d6: frame_vm_group_bin_2417 (RW)
0x1d7: frame_vm_group_bin_18507 (RW)
0x1d8: frame_vm_group_bin_11428 (RW)
0x1d9: frame_vm_group_bin_4244 (RW)
0x1d: frame_vm_group_bin_16649 (RW)
0x1da: frame_vm_group_bin_20343 (RW)
0x1db: frame_vm_group_bin_13146 (RW)
0x1dc: frame_vm_group_bin_4973 (RW)
0x1dd: frame_vm_group_bin_22154 (RW)
0x1de: frame_vm_group_bin_15005 (RW)
0x1df: frame_vm_group_bin_7789 (RW)
0x1e0: frame_vm_group_bin_0623 (RW)
0x1e1: frame_vm_group_bin_16820 (RW)
0x1e2: frame_vm_group_bin_9611 (RW)
0x1e3: frame_vm_group_bin_2450 (RW)
0x1e4: frame_vm_group_bin_18536 (RW)
0x1e5: frame_vm_group_bin_11462 (RW)
0x1e6: frame_vm_group_bin_4278 (RW)
0x1e7: frame_vm_group_bin_20376 (RW)
0x1e8: frame_vm_group_bin_13179 (RW)
0x1e9: frame_vm_group_bin_6022 (RW)
0x1e: frame_vm_group_bin_10318 (RW)
0x1ea: frame_vm_group_bin_22187 (RW)
0x1eb: frame_vm_group_bin_15036 (RW)
0x1ec: frame_vm_group_bin_7822 (RW)
0x1ed: frame_vm_group_bin_0657 (RW)
0x1ee: frame_vm_group_bin_16853 (RW)
0x1ef: frame_vm_group_bin_9644 (RW)
0x1f0: frame_vm_group_bin_2482 (RW)
0x1f1: frame_vm_group_bin_18561 (RW)
0x1f2: frame_vm_group_bin_11495 (RW)
0x1f3: frame_vm_group_bin_4311 (RW)
0x1f4: frame_vm_group_bin_20409 (RW)
0x1f5: frame_vm_group_bin_13212 (RW)
0x1f6: frame_vm_group_bin_14271 (RW)
0x1f7: frame_vm_group_bin_22220 (RW)
0x1f8: frame_vm_group_bin_15061 (RW)
0x1f9: frame_vm_group_bin_7854 (RW)
0x1f: frame_vm_group_bin_3158 (RW)
0x1fa: frame_vm_group_bin_0691 (RW)
0x1fb: frame_vm_group_bin_16886 (RW)
0x1fc: frame_vm_group_bin_9678 (RW)
0x1fd: frame_vm_group_bin_2516 (RW)
0x1fe: frame_vm_group_bin_18593 (RW)
0x1ff: frame_vm_group_bin_11529 (RW)
0x20: frame_vm_group_bin_19227 (RW)
0x21: frame_vm_group_bin_12055 (RW)
0x22: frame_vm_group_bin_4956 (RW)
0x23: frame_vm_group_bin_21053 (RW)
0x24: frame_vm_group_bin_13876 (RW)
0x25: frame_vm_group_bin_6695 (RW)
0x26: frame_vm_group_bin_22891 (RW)
0x27: frame_vm_group_bin_15708 (RW)
0x28: frame_vm_group_bin_8517 (RW)
0x29: frame_vm_group_bin_1325 (RW)
0x2: frame_vm_group_bin_1229 (RW)
0x2a: frame_vm_group_bin_17504 (RW)
0x2b: frame_vm_group_bin_10351 (RW)
0x2c: frame_vm_group_bin_3191 (RW)
0x2d: frame_vm_group_bin_19260 (RW)
0x2e: frame_vm_group_bin_12087 (RW)
0x2f: frame_vm_group_bin_4988 (RW)
0x30: frame_vm_group_bin_21086 (RW)
0x31: frame_vm_group_bin_13908 (RW)
0x32: frame_vm_group_bin_6727 (RW)
0x33: frame_vm_group_bin_22924 (RW)
0x34: frame_vm_group_bin_15741 (RW)
0x35: frame_vm_group_bin_8549 (RW)
0x36: frame_vm_group_bin_1358 (RW)
0x37: frame_vm_group_bin_17532 (RW)
0x38: frame_vm_group_bin_10383 (RW)
0x39: frame_vm_group_bin_3224 (RW)
0x3: frame_vm_group_bin_17440 (RW)
0x3a: frame_vm_group_bin_19294 (RW)
0x3b: frame_vm_group_bin_12120 (RW)
0x3c: frame_vm_group_bin_5022 (RW)
0x3d: frame_vm_group_bin_21120 (RW)
0x3e: frame_vm_group_bin_13942 (RW)
0x3f: frame_vm_group_bin_6760 (RW)
0x40: frame_vm_group_bin_22957 (RW)
0x41: frame_vm_group_bin_15775 (RW)
0x42: frame_vm_group_bin_8582 (RW)
0x43: frame_vm_group_bin_1393 (RW)
0x44: frame_vm_group_bin_7266 (RW)
0x45: frame_vm_group_bin_10411 (RW)
0x46: frame_vm_group_bin_3257 (RW)
0x47: frame_vm_group_bin_19327 (RW)
0x48: frame_vm_group_bin_12153 (RW)
0x49: frame_vm_group_bin_5055 (RW)
0x4: frame_vm_group_bin_10251 (RW)
0x4a: frame_vm_group_bin_21152 (RW)
0x4b: frame_vm_group_bin_13975 (RW)
0x4c: frame_vm_group_bin_6793 (RW)
0x4d: frame_vm_group_bin_22990 (RW)
0x4e: frame_vm_group_bin_15807 (RW)
0x4f: frame_vm_group_bin_8614 (RW)
0x50: frame_vm_group_bin_1426 (RW)
0x51: frame_vm_group_bin_11940 (RW)
0x52: frame_vm_group_bin_10439 (RW)
0x53: frame_vm_group_bin_3290 (RW)
0x54: frame_vm_group_bin_19360 (RW)
0x55: frame_vm_group_bin_12183 (RW)
0x56: frame_vm_group_bin_5089 (RW)
0x57: frame_vm_group_bin_21185 (RW)
0x58: frame_vm_group_bin_14008 (RW)
0x59: frame_vm_group_bin_6823 (RW)
0x5: frame_vm_group_bin_3092 (RW)
0x5a: frame_vm_group_bin_23023 (RW)
0x5b: frame_vm_group_bin_15840 (RW)
0x5c: frame_vm_group_bin_8648 (RW)
0x5d: frame_vm_group_bin_1460 (RW)
0x5e: frame_vm_group_bin_17602 (RW)
0x5f: frame_vm_group_bin_10471 (RW)
0x60: frame_vm_group_bin_3324 (RW)
0x61: frame_vm_group_bin_19394 (RW)
0x62: frame_vm_group_bin_12213 (RW)
0x63: frame_vm_group_bin_5123 (RW)
0x64: frame_vm_group_bin_21219 (RW)
0x65: frame_vm_group_bin_14042 (RW)
0x66: frame_vm_group_bin_6853 (RW)
0x67: frame_vm_group_bin_23056 (RW)
0x68: frame_vm_group_bin_15873 (RW)
0x69: frame_vm_group_bin_8682 (RW)
0x6: frame_vm_group_bin_19160 (RW)
0x6a: frame_vm_group_bin_1493 (RW)
0x6b: frame_vm_group_bin_17633 (RW)
0x6c: frame_vm_group_bin_10504 (RW)
0x6d: frame_vm_group_bin_3357 (RW)
0x6e: frame_vm_group_bin_19426 (RW)
0x6f: frame_vm_group_bin_12245 (RW)
0x70: frame_vm_group_bin_5156 (RW)
0x71: frame_vm_group_bin_21252 (RW)
0x72: frame_vm_group_bin_14075 (RW)
0x73: frame_vm_group_bin_6878 (RW)
0x74: frame_vm_group_bin_23089 (RW)
0x75: frame_vm_group_bin_15906 (RW)
0x76: frame_vm_group_bin_8715 (RW)
0x77: frame_vm_group_bin_1526 (RW)
0x78: frame_vm_group_bin_17666 (RW)
0x79: frame_vm_group_bin_10536 (RW)
0x7: frame_vm_group_bin_11996 (RW)
0x7a: frame_vm_group_bin_3388 (RW)
0x7b: frame_vm_group_bin_19457 (RW)
0x7c: frame_vm_group_bin_12279 (RW)
0x7d: frame_vm_group_bin_5190 (RW)
0x7e: frame_vm_group_bin_21286 (RW)
0x7f: frame_vm_group_bin_14109 (RW)
0x80: frame_vm_group_bin_6903 (RW)
0x81: frame_vm_group_bin_23123 (RW)
0x82: frame_vm_group_bin_15940 (RW)
0x83: frame_vm_group_bin_8749 (RW)
0x84: frame_vm_group_bin_1560 (RW)
0x85: frame_vm_group_bin_7290 (RW)
0x86: frame_vm_group_bin_10570 (RW)
0x87: frame_vm_group_bin_3415 (RW)
0x88: frame_vm_group_bin_19490 (RW)
0x89: frame_vm_group_bin_12312 (RW)
0x8: frame_vm_group_bin_4892 (RW)
0x8a: frame_vm_group_bin_5223 (RW)
0x8b: frame_vm_group_bin_21318 (RW)
0x8c: frame_vm_group_bin_14142 (RW)
0x8d: frame_vm_group_bin_6931 (RW)
0x8e: frame_vm_group_bin_23155 (RW)
0x8f: frame_vm_group_bin_15973 (RW)
0x90: frame_vm_group_bin_8782 (RW)
0x91: frame_vm_group_bin_1593 (RW)
0x92: frame_vm_group_bin_11963 (RW)
0x93: frame_vm_group_bin_10603 (RW)
0x94: frame_vm_group_bin_3437 (RW)
0x95: frame_vm_group_bin_19523 (RW)
0x96: frame_vm_group_bin_12344 (RW)
0x97: frame_vm_group_bin_5256 (RW)
0x98: frame_vm_group_bin_21350 (RW)
0x99: frame_vm_group_bin_14175 (RW)
0x9: frame_vm_group_bin_20985 (RW)
0x9a: frame_vm_group_bin_6963 (RW)
0x9b: frame_vm_group_bin_23188 (RW)
0x9c: frame_vm_group_bin_16009 (RW)
0x9d: frame_vm_group_bin_8816 (RW)
0x9e: frame_vm_group_bin_1627 (RW)
0x9f: frame_vm_group_bin_16695 (RW)
0xa0: frame_vm_group_bin_10637 (RW)
0xa1: frame_vm_group_bin_3463 (RW)
0xa2: frame_vm_group_bin_19557 (RW)
0xa3: frame_vm_group_bin_12378 (RW)
0xa4: frame_vm_group_bin_5290 (RW)
0xa5: frame_vm_group_bin_21384 (RW)
0xa6: frame_vm_group_bin_14208 (RW)
0xa7: frame_vm_group_bin_6995 (RW)
0xa8: frame_vm_group_bin_23215 (RW)
0xa9: frame_vm_group_bin_16042 (RW)
0xa: frame_vm_group_bin_13816 (RW)
0xaa: frame_vm_group_bin_8849 (RW)
0xab: frame_vm_group_bin_1660 (RW)
0xac: frame_vm_group_bin_21329 (RW)
0xad: frame_vm_group_bin_10668 (RW)
0xae: frame_vm_group_bin_3489 (RW)
0xaf: frame_vm_group_bin_19591 (RW)
0xb0: frame_vm_group_bin_12411 (RW)
0xb1: frame_vm_group_bin_5322 (RW)
0xb2: frame_vm_group_bin_21417 (RW)
0xb3: frame_vm_group_bin_14241 (RW)
0xb4: frame_vm_group_bin_7028 (RW)
0xb5: frame_vm_group_bin_23237 (RW)
0xb6: frame_vm_group_bin_16075 (RW)
0xb7: frame_vm_group_bin_8881 (RW)
0xb8: frame_vm_group_bin_1693 (RW)
0xb9: frame_vm_group_bin_2704 (RW)
0xb: frame_vm_group_bin_6628 (RW)
0xba: frame_vm_group_bin_10702 (RW)
0xbb: frame_vm_group_bin_3517 (RW)
0xbc: frame_vm_group_bin_19625 (RW)
0xbd: frame_vm_group_bin_12444 (RW)
0xbe: frame_vm_group_bin_5354 (RW)
0xbf: frame_vm_group_bin_21450 (RW)
0xc0: frame_vm_group_bin_14274 (RW)
0xc1: frame_vm_group_bin_7060 (RW)
0xc2: frame_vm_group_bin_1361 (RW)
0xc3: frame_vm_group_bin_16108 (RW)
0xc4: frame_vm_group_bin_8914 (RW)
0xc5: frame_vm_group_bin_1726 (RW)
0xc6: frame_vm_group_bin_7314 (RW)
0xc7: frame_vm_group_bin_10734 (RW)
0xc8: frame_vm_group_bin_3548 (RW)
0xc9: frame_vm_group_bin_19655 (RW)
0xc: frame_vm_group_bin_22824 (RW)
0xca: frame_vm_group_bin_12476 (RW)
0xcb: frame_vm_group_bin_5386 (RW)
0xcc: frame_vm_group_bin_21482 (RW)
0xcd: frame_vm_group_bin_14305 (RW)
0xce: frame_vm_group_bin_7092 (RW)
0xcf: frame_vm_group_bin_17727 (RW)
0xd0: frame_vm_group_bin_16139 (RW)
0xd1: frame_vm_group_bin_8946 (RW)
0xd2: frame_vm_group_bin_1758 (RW)
0xd3: frame_vm_group_bin_11987 (RW)
0xd4: frame_vm_group_bin_10767 (RW)
0xd5: frame_vm_group_bin_3580 (RW)
0xd6: frame_vm_group_bin_19682 (RW)
0xd7: frame_vm_group_bin_12509 (RW)
0xd8: frame_vm_group_bin_5419 (RW)
0xd9: frame_vm_group_bin_21514 (RW)
0xd: frame_vm_group_bin_15641 (RW)
0xda: frame_vm_group_bin_14339 (RW)
0xdb: frame_vm_group_bin_7125 (RW)
0xdc: frame_vm_group_bin_22432 (RW)
0xdd: frame_vm_group_bin_16173 (RW)
0xde: frame_vm_group_bin_8980 (RW)
0xdf: frame_vm_group_bin_1792 (RW)
0xe0: frame_vm_group_bin_17895 (RW)
0xe1: frame_vm_group_bin_10800 (RW)
0xe2: frame_vm_group_bin_3615 (RW)
0xe3: frame_vm_group_bin_19715 (RW)
0xe4: frame_vm_group_bin_12543 (RW)
0xe5: frame_vm_group_bin_5452 (RW)
0xe6: frame_vm_group_bin_21548 (RW)
0xe7: frame_vm_group_bin_14372 (RW)
0xe8: frame_vm_group_bin_7157 (RW)
0xe9: frame_vm_group_bin_3797 (RW)
0xe: frame_vm_group_bin_8451 (RW)
0xea: frame_vm_group_bin_16204 (RW)
0xeb: frame_vm_group_bin_9013 (RW)
0xec: frame_vm_group_bin_1825 (RW)
0xed: frame_vm_group_bin_17927 (RW)
0xee: frame_vm_group_bin_10833 (RW)
0xef: frame_vm_group_bin_3648 (RW)
0xf0: frame_vm_group_bin_19748 (RW)
0xf1: frame_vm_group_bin_12576 (RW)
0xf2: frame_vm_group_bin_5484 (RW)
0xf3: frame_vm_group_bin_21581 (RW)
0xf4: frame_vm_group_bin_14405 (RW)
0xf5: frame_vm_group_bin_7192 (RW)
0xf6: frame_vm_group_bin_8437 (RW)
0xf7: frame_vm_group_bin_16231 (RW)
0xf8: frame_vm_group_bin_9046 (RW)
0xf9: frame_vm_group_bin_1858 (RW)
0xf: frame_vm_group_bin_1261 (RW)
0xfa: frame_vm_group_bin_17959 (RW)
0xfb: frame_vm_group_bin_10867 (RW)
0xfc: frame_vm_group_bin_3682 (RW)
0xfd: frame_vm_group_bin_19782 (RW)
0xfe: frame_vm_group_bin_12610 (RW)
0xff: frame_vm_group_bin_5517 (RW)
}
pt_vm_group_bin_0272 {
0x0: frame_vm_group_bin_14887 (RW)
0x100: frame_vm_group_bin_20879 (RW)
0x101: frame_vm_group_bin_13692 (RW)
0x102: frame_vm_group_bin_6503 (RW)
0x103: frame_vm_group_bin_22700 (RW)
0x104: frame_vm_group_bin_15517 (RW)
0x105: frame_vm_group_bin_8326 (RW)
0x106: frame_vm_group_bin_1137 (RW)
0x107: frame_vm_group_bin_17362 (RW)
0x108: frame_vm_group_bin_10159 (RW)
0x109: frame_vm_group_bin_3000 (RW)
0x10: frame_vm_group_bin_16735 (RW)
0x10a: frame_vm_group_bin_19070 (RW)
0x10b: frame_vm_group_bin_1625 (RW)
0x10c: frame_vm_group_bin_4801 (RW)
0x10d: frame_vm_group_bin_20906 (RW)
0x10e: frame_vm_group_bin_13724 (RW)
0x10f: frame_vm_group_bin_6536 (RW)
0x110: frame_vm_group_bin_22733 (RW)
0x111: frame_vm_group_bin_15549 (RW)
0x112: frame_vm_group_bin_8359 (RW)
0x113: frame_vm_group_bin_1170 (RW)
0x114: frame_vm_group_bin_17392 (RW)
0x115: frame_vm_group_bin_10192 (RW)
0x116: frame_vm_group_bin_3033 (RW)
0x117: frame_vm_group_bin_19103 (RW)
0x118: frame_vm_group_bin_6265 (RW)
0x119: frame_vm_group_bin_4833 (RW)
0x11: frame_vm_group_bin_9526 (RW)
0x11a: frame_vm_group_bin_20935 (RW)
0x11b: frame_vm_group_bin_13759 (RW)
0x11c: frame_vm_group_bin_6570 (RW)
0x11d: frame_vm_group_bin_22766 (RW)
0x11e: frame_vm_group_bin_15583 (RW)
0x11f: frame_vm_group_bin_8393 (RW)
0x120: frame_vm_group_bin_1204 (RW)
0x121: frame_vm_group_bin_17420 (RW)
0x122: frame_vm_group_bin_10226 (RW)
0x123: frame_vm_group_bin_3067 (RW)
0x124: frame_vm_group_bin_19135 (RW)
0x125: frame_vm_group_bin_11972 (RW)
0x126: frame_vm_group_bin_4867 (RW)
0x127: frame_vm_group_bin_20962 (RW)
0x128: frame_vm_group_bin_13792 (RW)
0x129: frame_vm_group_bin_6603 (RW)
0x12: frame_vm_group_bin_2366 (RW)
0x12a: frame_vm_group_bin_22799 (RW)
0x12b: frame_vm_group_bin_15616 (RW)
0x12c: frame_vm_group_bin_8426 (RW)
0x12d: frame_vm_group_bin_1237 (RW)
0x12e: frame_vm_group_bin_17445 (RW)
0x12f: frame_vm_group_bin_10259 (RW)
0x130: frame_vm_group_bin_3100 (RW)
0x131: frame_vm_group_bin_19168 (RW)
0x132: frame_vm_group_bin_12004 (RW)
0x133: frame_vm_group_bin_4900 (RW)
0x134: frame_vm_group_bin_20993 (RW)
0x135: frame_vm_group_bin_13823 (RW)
0x136: frame_vm_group_bin_6636 (RW)
0x137: frame_vm_group_bin_22832 (RW)
0x138: frame_vm_group_bin_15649 (RW)
0x139: frame_vm_group_bin_8459 (RW)
0x13: frame_vm_group_bin_18465 (RW)
0x13a: frame_vm_group_bin_1270 (RW)
0x13b: frame_vm_group_bin_2751 (RW)
0x13c: frame_vm_group_bin_10293 (RW)
0x13d: frame_vm_group_bin_3133 (RW)
0x13e: frame_vm_group_bin_19202 (RW)
0x13f: frame_vm_group_bin_12035 (RW)
0x140: frame_vm_group_bin_4932 (RW)
0x141: frame_vm_group_bin_21027 (RW)
0x142: frame_vm_group_bin_13854 (RW)
0x143: frame_vm_group_bin_6670 (RW)
0x144: frame_vm_group_bin_22866 (RW)
0x145: frame_vm_group_bin_15683 (RW)
0x146: frame_vm_group_bin_8493 (RW)
0x147: frame_vm_group_bin_1301 (RW)
0x148: frame_vm_group_bin_7362 (RW)
0x149: frame_vm_group_bin_10326 (RW)
0x14: frame_vm_group_bin_6182 (RW)
0x14a: frame_vm_group_bin_3166 (RW)
0x14b: frame_vm_group_bin_19235 (RW)
0x14c: frame_vm_group_bin_12062 (RW)
0x14d: frame_vm_group_bin_0231 (RW)
0x14e: frame_vm_group_bin_21061 (RW)
0x14f: frame_vm_group_bin_13883 (RW)
0x150: frame_vm_group_bin_6703 (RW)
0x151: frame_vm_group_bin_22899 (RW)
0x152: frame_vm_group_bin_15716 (RW)
0x153: frame_vm_group_bin_8525 (RW)
0x154: frame_vm_group_bin_1333 (RW)
0x155: frame_vm_group_bin_17512 (RW)
0x156: frame_vm_group_bin_10359 (RW)
0x157: frame_vm_group_bin_3199 (RW)
0x158: frame_vm_group_bin_19268 (RW)
0x159: frame_vm_group_bin_12095 (RW)
0x15: frame_vm_group_bin_4194 (RW)
0x15a: frame_vm_group_bin_4997 (RW)
0x15b: frame_vm_group_bin_21095 (RW)
0x15c: frame_vm_group_bin_13917 (RW)
0x15d: frame_vm_group_bin_6736 (RW)
0x15e: frame_vm_group_bin_22933 (RW)
0x15f: frame_vm_group_bin_15750 (RW)
0x160: frame_vm_group_bin_8557 (RW)
0x161: frame_vm_group_bin_1368 (RW)
0x162: frame_vm_group_bin_16767 (RW)
0x163: frame_vm_group_bin_10392 (RW)
0x164: frame_vm_group_bin_3232 (RW)
0x165: frame_vm_group_bin_19302 (RW)
0x166: frame_vm_group_bin_12128 (RW)
0x167: frame_vm_group_bin_5030 (RW)
0x168: frame_vm_group_bin_21128 (RW)
0x169: frame_vm_group_bin_13950 (RW)
0x16: frame_vm_group_bin_20289 (RW)
0x16a: frame_vm_group_bin_6768 (RW)
0x16b: frame_vm_group_bin_22965 (RW)
0x16c: frame_vm_group_bin_15783 (RW)
0x16d: frame_vm_group_bin_8590 (RW)
0x16e: frame_vm_group_bin_1401 (RW)
0x16f: frame_vm_group_bin_21399 (RW)
0x170: frame_vm_group_bin_10417 (RW)
0x171: frame_vm_group_bin_3265 (RW)
0x172: frame_vm_group_bin_19335 (RW)
0x173: frame_vm_group_bin_12160 (RW)
0x174: frame_vm_group_bin_5063 (RW)
0x175: frame_vm_group_bin_21160 (RW)
0x176: frame_vm_group_bin_13983 (RW)
0x177: frame_vm_group_bin_6801 (RW)
0x178: frame_vm_group_bin_22998 (RW)
0x179: frame_vm_group_bin_15815 (RW)
0x17: frame_vm_group_bin_13094 (RW)
0x17a: frame_vm_group_bin_8623 (RW)
0x17b: frame_vm_group_bin_1435 (RW)
0x17c: frame_vm_group_bin_17586 (RW)
0x17d: frame_vm_group_bin_10446 (RW)
0x17e: frame_vm_group_bin_3299 (RW)
0x17f: frame_vm_group_bin_19369 (RW)
0x180: frame_vm_group_bin_12191 (RW)
0x181: frame_vm_group_bin_5098 (RW)
0x182: frame_vm_group_bin_21194 (RW)
0x183: frame_vm_group_bin_14017 (RW)
0x184: frame_vm_group_bin_6832 (RW)
0x185: frame_vm_group_bin_23031 (RW)
0x186: frame_vm_group_bin_15848 (RW)
0x187: frame_vm_group_bin_8656 (RW)
0x188: frame_vm_group_bin_1468 (RW)
0x189: frame_vm_group_bin_17609 (RW)
0x18: frame_vm_group_bin_0460 (RW)
0x18a: frame_vm_group_bin_10479 (RW)
0x18b: frame_vm_group_bin_3332 (RW)
0x18c: frame_vm_group_bin_19402 (RW)
0x18d: frame_vm_group_bin_12221 (RW)
0x18e: frame_vm_group_bin_5131 (RW)
0x18f: frame_vm_group_bin_21227 (RW)
0x190: frame_vm_group_bin_14050 (RW)
0x191: frame_vm_group_bin_6859 (RW)
0x192: frame_vm_group_bin_23064 (RW)
0x193: frame_vm_group_bin_15881 (RW)
0x194: frame_vm_group_bin_8690 (RW)
0x195: frame_vm_group_bin_1501 (RW)
0x196: frame_vm_group_bin_17641 (RW)
0x197: frame_vm_group_bin_10512 (RW)
0x198: frame_vm_group_bin_3365 (RW)
0x199: frame_vm_group_bin_19434 (RW)
0x19: frame_vm_group_bin_22102 (RW)
0x19a: frame_vm_group_bin_12254 (RW)
0x19b: frame_vm_group_bin_5165 (RW)
0x19c: frame_vm_group_bin_21261 (RW)
0x19d: frame_vm_group_bin_14084 (RW)
0x19e: frame_vm_group_bin_6885 (RW)
0x19f: frame_vm_group_bin_23098 (RW)
0x1: frame_vm_group_bin_7672 (RW)
0x1a0: frame_vm_group_bin_15915 (RW)
0x1a1: frame_vm_group_bin_8724 (RW)
0x1a2: frame_vm_group_bin_1535 (RW)
0x1a3: frame_vm_group_bin_17675 (RW)
0x1a4: frame_vm_group_bin_10545 (RW)
0x1a5: frame_vm_group_bin_3396 (RW)
0x1a6: frame_vm_group_bin_19465 (RW)
0x1a7: frame_vm_group_bin_12287 (RW)
0x1a8: frame_vm_group_bin_5198 (RW)
0x1a9: frame_vm_group_bin_21294 (RW)
0x1a: frame_vm_group_bin_14954 (RW)
0x1aa: frame_vm_group_bin_14117 (RW)
0x1ab: frame_vm_group_bin_6908 (RW)
0x1ac: frame_vm_group_bin_23131 (RW)
0x1ad: frame_vm_group_bin_15948 (RW)
0x1ae: frame_vm_group_bin_8757 (RW)
0x1af: frame_vm_group_bin_1568 (RW)
0x1b0: frame_vm_group_bin_21423 (RW)
0x1b1: frame_vm_group_bin_10578 (RW)
0x1b2: frame_vm_group_bin_3420 (RW)
0x1b3: frame_vm_group_bin_19498 (RW)
0x1b4: frame_vm_group_bin_12320 (RW)
0x1b5: frame_vm_group_bin_5231 (RW)
0x1b6: frame_vm_group_bin_21326 (RW)
0x1b7: frame_vm_group_bin_14150 (RW)
0x1b8: frame_vm_group_bin_6938 (RW)
0x1b9: frame_vm_group_bin_23163 (RW)
0x1b: frame_vm_group_bin_7738 (RW)
0x1ba: frame_vm_group_bin_15984 (RW)
0x1bb: frame_vm_group_bin_8791 (RW)
0x1bc: frame_vm_group_bin_1602 (RW)
0x1bd: frame_vm_group_bin_17729 (RW)
0x1be: frame_vm_group_bin_10612 (RW)
0x1bf: frame_vm_group_bin_3443 (RW)
0x1c0: frame_vm_group_bin_19532 (RW)
0x1c1: frame_vm_group_bin_12353 (RW)
0x1c2: frame_vm_group_bin_5265 (RW)
0x1c3: frame_vm_group_bin_21359 (RW)
0x1c4: frame_vm_group_bin_14183 (RW)
0x1c5: frame_vm_group_bin_6970 (RW)
0x1c6: frame_vm_group_bin_23196 (RW)
0x1c7: frame_vm_group_bin_16017 (RW)
0x1c8: frame_vm_group_bin_8824 (RW)
0x1c9: frame_vm_group_bin_1635 (RW)
0x1c: frame_vm_group_bin_0575 (RW)
0x1ca: frame_vm_group_bin_17756 (RW)
0x1cb: frame_vm_group_bin_5990 (RW)
0x1cc: frame_vm_group_bin_3468 (RW)
0x1cd: frame_vm_group_bin_19565 (RW)
0x1ce: frame_vm_group_bin_12386 (RW)
0x1cf: frame_vm_group_bin_5298 (RW)
0x1d0: frame_vm_group_bin_21392 (RW)
0x1d1: frame_vm_group_bin_14216 (RW)
0x1d2: frame_vm_group_bin_7003 (RW)
0x1d3: frame_vm_group_bin_23220 (RW)
0x1d4: frame_vm_group_bin_16050 (RW)
0x1d5: frame_vm_group_bin_8857 (RW)
0x1d6: frame_vm_group_bin_1668 (RW)
0x1d7: frame_vm_group_bin_17786 (RW)
0x1d8: frame_vm_group_bin_10676 (RW)
0x1d9: frame_vm_group_bin_3494 (RW)
0x1d: frame_vm_group_bin_16769 (RW)
0x1da: frame_vm_group_bin_19600 (RW)
0x1db: frame_vm_group_bin_12420 (RW)
0x1dc: frame_vm_group_bin_5330 (RW)
0x1dd: frame_vm_group_bin_21425 (RW)
0x1de: frame_vm_group_bin_14249 (RW)
0x1df: frame_vm_group_bin_7036 (RW)
0x1e0: frame_vm_group_bin_23242 (RW)
0x1e1: frame_vm_group_bin_16083 (RW)
0x1e2: frame_vm_group_bin_8889 (RW)
0x1e3: frame_vm_group_bin_1701 (RW)
0x1e4: frame_vm_group_bin_17816 (RW)
0x1e5: frame_vm_group_bin_10709 (RW)
0x1e6: frame_vm_group_bin_3523 (RW)
0x1e7: frame_vm_group_bin_19632 (RW)
0x1e8: frame_vm_group_bin_12451 (RW)
0x1e9: frame_vm_group_bin_5361 (RW)
0x1e: frame_vm_group_bin_9560 (RW)
0x1ea: frame_vm_group_bin_21457 (RW)
0x1eb: frame_vm_group_bin_14281 (RW)
0x1ec: frame_vm_group_bin_7067 (RW)
0x1ed: frame_vm_group_bin_3893 (RW)
0x1ee: frame_vm_group_bin_16115 (RW)
0x1ef: frame_vm_group_bin_8921 (RW)
0x1f0: frame_vm_group_bin_1733 (RW)
0x1f1: frame_vm_group_bin_21448 (RW)
0x1f2: frame_vm_group_bin_10741 (RW)
0x1f3: frame_vm_group_bin_3555 (RW)
0x1f4: frame_vm_group_bin_19660 (RW)
0x1f5: frame_vm_group_bin_12483 (RW)
0x1f6: frame_vm_group_bin_5393 (RW)
0x1f7: frame_vm_group_bin_21489 (RW)
0x1f8: frame_vm_group_bin_14312 (RW)
0x1f9: frame_vm_group_bin_7099 (RW)
0x1f: frame_vm_group_bin_2400 (RW)
0x1fa: frame_vm_group_bin_8532 (RW)
0x1fb: frame_vm_group_bin_16147 (RW)
0x1fc: frame_vm_group_bin_8954 (RW)
0x1fd: frame_vm_group_bin_1766 (RW)
0x1fe: frame_vm_group_bin_2822 (RW)
0x1ff: frame_vm_group_bin_10774 (RW)
0x20: frame_vm_group_bin_18494 (RW)
0x21: frame_vm_group_bin_11411 (RW)
0x22: frame_vm_group_bin_4227 (RW)
0x23: frame_vm_group_bin_20325 (RW)
0x24: frame_vm_group_bin_13128 (RW)
0x25: frame_vm_group_bin_5975 (RW)
0x26: frame_vm_group_bin_22136 (RW)
0x27: frame_vm_group_bin_14987 (RW)
0x28: frame_vm_group_bin_7771 (RW)
0x29: frame_vm_group_bin_0607 (RW)
0x2: frame_vm_group_bin_0511 (RW)
0x2a: frame_vm_group_bin_16802 (RW)
0x2b: frame_vm_group_bin_9593 (RW)
0x2c: frame_vm_group_bin_2432 (RW)
0x2d: frame_vm_group_bin_18521 (RW)
0x2e: frame_vm_group_bin_11444 (RW)
0x2f: frame_vm_group_bin_4260 (RW)
0x30: frame_vm_group_bin_20358 (RW)
0x31: frame_vm_group_bin_13161 (RW)
0x32: frame_vm_group_bin_6006 (RW)
0x33: frame_vm_group_bin_22169 (RW)
0x34: frame_vm_group_bin_15020 (RW)
0x35: frame_vm_group_bin_7804 (RW)
0x36: frame_vm_group_bin_0638 (RW)
0x37: frame_vm_group_bin_16835 (RW)
0x38: frame_vm_group_bin_9626 (RW)
0x39: frame_vm_group_bin_2465 (RW)
0x3: frame_vm_group_bin_16701 (RW)
0x3a: frame_vm_group_bin_18546 (RW)
0x3b: frame_vm_group_bin_11478 (RW)
0x3c: frame_vm_group_bin_4294 (RW)
0x3d: frame_vm_group_bin_20392 (RW)
0x3e: frame_vm_group_bin_13195 (RW)
0x3f: frame_vm_group_bin_6038 (RW)
0x40: frame_vm_group_bin_22203 (RW)
0x41: frame_vm_group_bin_15049 (RW)
0x42: frame_vm_group_bin_7837 (RW)
0x43: frame_vm_group_bin_0673 (RW)
0x44: frame_vm_group_bin_16868 (RW)
0x45: frame_vm_group_bin_9660 (RW)
0x46: frame_vm_group_bin_2498 (RW)
0x47: frame_vm_group_bin_18575 (RW)
0x48: frame_vm_group_bin_11511 (RW)
0x49: frame_vm_group_bin_4327 (RW)
0x4: frame_vm_group_bin_9493 (RW)
0x4a: frame_vm_group_bin_20425 (RW)
0x4b: frame_vm_group_bin_13228 (RW)
0x4c: frame_vm_group_bin_19106 (RW)
0x4d: frame_vm_group_bin_22236 (RW)
0x4e: frame_vm_group_bin_15073 (RW)
0x4f: frame_vm_group_bin_7870 (RW)
0x50: frame_vm_group_bin_0706 (RW)
0x51: frame_vm_group_bin_16900 (RW)
0x52: frame_vm_group_bin_9692 (RW)
0x53: frame_vm_group_bin_2531 (RW)
0x54: frame_vm_group_bin_18608 (RW)
0x55: frame_vm_group_bin_11544 (RW)
0x56: frame_vm_group_bin_4362 (RW)
0x57: frame_vm_group_bin_20458 (RW)
0x58: frame_vm_group_bin_13261 (RW)
0x59: frame_vm_group_bin_0483 (RW)
0x5: frame_vm_group_bin_2333 (RW)
0x5a: frame_vm_group_bin_22270 (RW)
0x5b: frame_vm_group_bin_15098 (RW)
0x5c: frame_vm_group_bin_7904 (RW)
0x5d: frame_vm_group_bin_0740 (RW)
0x5e: frame_vm_group_bin_16934 (RW)
0x5f: frame_vm_group_bin_9726 (RW)
0x60: frame_vm_group_bin_2565 (RW)
0x61: frame_vm_group_bin_18641 (RW)
0x62: frame_vm_group_bin_11575 (RW)
0x63: frame_vm_group_bin_4396 (RW)
0x64: frame_vm_group_bin_20492 (RW)
0x65: frame_vm_group_bin_13295 (RW)
0x66: frame_vm_group_bin_6120 (RW)
0x67: frame_vm_group_bin_22302 (RW)
0x68: frame_vm_group_bin_15127 (RW)
0x69: frame_vm_group_bin_7938 (RW)
0x6: frame_vm_group_bin_18434 (RW)
0x6a: frame_vm_group_bin_0773 (RW)
0x6b: frame_vm_group_bin_16967 (RW)
0x6c: frame_vm_group_bin_9759 (RW)
0x6d: frame_vm_group_bin_2598 (RW)
0x6e: frame_vm_group_bin_18674 (RW)
0x6f: frame_vm_group_bin_11600 (RW)
0x70: frame_vm_group_bin_4429 (RW)
0x71: frame_vm_group_bin_20525 (RW)
0x72: frame_vm_group_bin_13327 (RW)
0x73: frame_vm_group_bin_6152 (RW)
0x74: frame_vm_group_bin_22335 (RW)
0x75: frame_vm_group_bin_15150 (RW)
0x76: frame_vm_group_bin_7971 (RW)
0x77: frame_vm_group_bin_0806 (RW)
0x78: frame_vm_group_bin_17000 (RW)
0x79: frame_vm_group_bin_9792 (RW)
0x7: frame_vm_group_bin_11346 (RW)
0x7a: frame_vm_group_bin_2632 (RW)
0x7b: frame_vm_group_bin_18707 (RW)
0x7c: frame_vm_group_bin_20315 (RW)
0x7d: frame_vm_group_bin_4463 (RW)
0x7e: frame_vm_group_bin_20559 (RW)
0x7f: frame_vm_group_bin_13361 (RW)
0x80: frame_vm_group_bin_6185 (RW)
0x81: frame_vm_group_bin_22368 (RW)
0x82: frame_vm_group_bin_15184 (RW)
0x83: frame_vm_group_bin_8003 (RW)
0x84: frame_vm_group_bin_0839 (RW)
0x85: frame_vm_group_bin_17034 (RW)
0x86: frame_vm_group_bin_9826 (RW)
0x87: frame_vm_group_bin_2665 (RW)
0x88: frame_vm_group_bin_18738 (RW)
0x89: frame_vm_group_bin_1576 (RW)
0x8: frame_vm_group_bin_4161 (RW)
0x8a: frame_vm_group_bin_4496 (RW)
0x8b: frame_vm_group_bin_20592 (RW)
0x8c: frame_vm_group_bin_13392 (RW)
0x8d: frame_vm_group_bin_19128 (RW)
0x8e: frame_vm_group_bin_22401 (RW)
0x8f: frame_vm_group_bin_15217 (RW)
0x90: frame_vm_group_bin_8031 (RW)
0x91: frame_vm_group_bin_0872 (RW)
0x92: frame_vm_group_bin_17067 (RW)
0x93: frame_vm_group_bin_9859 (RW)
0x94: frame_vm_group_bin_2698 (RW)
0x95: frame_vm_group_bin_18771 (RW)
0x96: frame_vm_group_bin_6221 (RW)
0x97: frame_vm_group_bin_4529 (RW)
0x98: frame_vm_group_bin_20625 (RW)
0x99: frame_vm_group_bin_13425 (RW)
0x9: frame_vm_group_bin_20257 (RW)
0x9a: frame_vm_group_bin_6243 (RW)
0x9b: frame_vm_group_bin_22434 (RW)
0x9c: frame_vm_group_bin_15252 (RW)
0x9d: frame_vm_group_bin_8062 (RW)
0x9e: frame_vm_group_bin_0906 (RW)
0x9f: frame_vm_group_bin_17101 (RW)
0xa0: frame_vm_group_bin_9892 (RW)
0xa1: frame_vm_group_bin_2732 (RW)
0xa2: frame_vm_group_bin_18805 (RW)
0xa3: frame_vm_group_bin_10961 (RW)
0xa4: frame_vm_group_bin_4562 (RW)
0xa5: frame_vm_group_bin_20658 (RW)
0xa6: frame_vm_group_bin_13459 (RW)
0xa7: frame_vm_group_bin_6274 (RW)
0xa8: frame_vm_group_bin_22467 (RW)
0xa9: frame_vm_group_bin_15284 (RW)
0xa: frame_vm_group_bin_13061 (RW)
0xaa: frame_vm_group_bin_8094 (RW)
0xab: frame_vm_group_bin_0939 (RW)
0xac: frame_vm_group_bin_17134 (RW)
0xad: frame_vm_group_bin_9925 (RW)
0xae: frame_vm_group_bin_2765 (RW)
0xaf: frame_vm_group_bin_18839 (RW)
0xb0: frame_vm_group_bin_15605 (RW)
0xb1: frame_vm_group_bin_4587 (RW)
0xb2: frame_vm_group_bin_20691 (RW)
0xb3: frame_vm_group_bin_13492 (RW)
0xb4: frame_vm_group_bin_6307 (RW)
0xb5: frame_vm_group_bin_22500 (RW)
0xb6: frame_vm_group_bin_15317 (RW)
0xb7: frame_vm_group_bin_8126 (RW)
0xb8: frame_vm_group_bin_0972 (RW)
0xb9: frame_vm_group_bin_17166 (RW)
0xb: frame_vm_group_bin_19083 (RW)
0xba: frame_vm_group_bin_9957 (RW)
0xbb: frame_vm_group_bin_2799 (RW)
0xbc: frame_vm_group_bin_18873 (RW)
0xbd: frame_vm_group_bin_20247 (RW)
0xbe: frame_vm_group_bin_4611 (RW)
0xbf: frame_vm_group_bin_20725 (RW)
0xc0: frame_vm_group_bin_13526 (RW)
0xc1: frame_vm_group_bin_6340 (RW)
0xc2: frame_vm_group_bin_22533 (RW)
0xc3: frame_vm_group_bin_15351 (RW)
0xc4: frame_vm_group_bin_8160 (RW)
0xc5: frame_vm_group_bin_1006 (RW)
0xc6: frame_vm_group_bin_17197 (RW)
0xc7: frame_vm_group_bin_9990 (RW)
0xc8: frame_vm_group_bin_2832 (RW)
0xc9: frame_vm_group_bin_18906 (RW)
0xc: frame_vm_group_bin_22072 (RW)
0xca: frame_vm_group_bin_1600 (RW)
0xcb: frame_vm_group_bin_4637 (RW)
0xcc: frame_vm_group_bin_20758 (RW)
0xcd: frame_vm_group_bin_13559 (RW)
0xce: frame_vm_group_bin_6372 (RW)
0xcf: frame_vm_group_bin_22566 (RW)
0xd0: frame_vm_group_bin_15384 (RW)
0xd1: frame_vm_group_bin_8193 (RW)
0xd2: frame_vm_group_bin_1031 (RW)
0xd3: frame_vm_group_bin_17230 (RW)
0xd4: frame_vm_group_bin_10023 (RW)
0xd5: frame_vm_group_bin_2864 (RW)
0xd6: frame_vm_group_bin_18939 (RW)
0xd7: frame_vm_group_bin_11796 (RW)
0xd8: frame_vm_group_bin_4670 (RW)
0xd9: frame_vm_group_bin_20791 (RW)
0xd: frame_vm_group_bin_14920 (RW)
0xda: frame_vm_group_bin_13593 (RW)
0xdb: frame_vm_group_bin_6404 (RW)
0xdc: frame_vm_group_bin_22600 (RW)
0xdd: frame_vm_group_bin_15418 (RW)
0xde: frame_vm_group_bin_8227 (RW)
0xdf: frame_vm_group_bin_1054 (RW)
0xe0: frame_vm_group_bin_17263 (RW)
0xe1: frame_vm_group_bin_10057 (RW)
0xe2: frame_vm_group_bin_2900 (RW)
0xe3: frame_vm_group_bin_18970 (RW)
0xe4: frame_vm_group_bin_11829 (RW)
0xe5: frame_vm_group_bin_4702 (RW)
0xe6: frame_vm_group_bin_20824 (RW)
0xe7: frame_vm_group_bin_13626 (RW)
0xe8: frame_vm_group_bin_6436 (RW)
0xe9: frame_vm_group_bin_22633 (RW)
0xe: frame_vm_group_bin_7705 (RW)
0xea: frame_vm_group_bin_15451 (RW)
0xeb: frame_vm_group_bin_8260 (RW)
0xec: frame_vm_group_bin_1077 (RW)
0xed: frame_vm_group_bin_17296 (RW)
0xee: frame_vm_group_bin_10090 (RW)
0xef: frame_vm_group_bin_2933 (RW)
0xf0: frame_vm_group_bin_19003 (RW)
0xf1: frame_vm_group_bin_11858 (RW)
0xf2: frame_vm_group_bin_4734 (RW)
0xf3: frame_vm_group_bin_20853 (RW)
0xf4: frame_vm_group_bin_13658 (RW)
0xf5: frame_vm_group_bin_6469 (RW)
0xf6: frame_vm_group_bin_22666 (RW)
0xf7: frame_vm_group_bin_15484 (RW)
0xf8: frame_vm_group_bin_8292 (RW)
0xf9: frame_vm_group_bin_1104 (RW)
0xf: frame_vm_group_bin_0543 (RW)
0xfa: frame_vm_group_bin_17330 (RW)
0xfb: frame_vm_group_bin_10124 (RW)
0xfc: frame_vm_group_bin_2967 (RW)
0xfd: frame_vm_group_bin_19037 (RW)
0xfe: frame_vm_group_bin_20270 (RW)
0xff: frame_vm_group_bin_4768 (RW)
}
pt_vm_group_bin_0328 {
0x0: frame_vm_group_bin_0286 (RW)
0x100: frame_vm_group_bin_6270 (RW)
0x101: frame_vm_group_bin_22463 (RW)
0x102: frame_vm_group_bin_15280 (RW)
0x103: frame_vm_group_bin_8090 (RW)
0x104: frame_vm_group_bin_0935 (RW)
0x105: frame_vm_group_bin_17130 (RW)
0x106: frame_vm_group_bin_9921 (RW)
0x107: frame_vm_group_bin_2761 (RW)
0x108: frame_vm_group_bin_18835 (RW)
0x109: frame_vm_group_bin_11721 (RW)
0x10: frame_vm_group_bin_2137 (RW)
0x10a: frame_vm_group_bin_3107 (RW)
0x10b: frame_vm_group_bin_20687 (RW)
0x10c: frame_vm_group_bin_13488 (RW)
0x10d: frame_vm_group_bin_6303 (RW)
0x10e: frame_vm_group_bin_22496 (RW)
0x10f: frame_vm_group_bin_15313 (RW)
0x110: frame_vm_group_bin_8122 (RW)
0x111: frame_vm_group_bin_0968 (RW)
0x112: frame_vm_group_bin_17162 (RW)
0x113: frame_vm_group_bin_9952 (RW)
0x114: frame_vm_group_bin_2794 (RW)
0x115: frame_vm_group_bin_18868 (RW)
0x116: frame_vm_group_bin_11743 (RW)
0x117: frame_vm_group_bin_4606 (RW)
0x118: frame_vm_group_bin_20720 (RW)
0x119: frame_vm_group_bin_13521 (RW)
0x11: frame_vm_group_bin_18231 (RW)
0x11a: frame_vm_group_bin_6336 (RW)
0x11b: frame_vm_group_bin_22529 (RW)
0x11c: frame_vm_group_bin_15347 (RW)
0x11d: frame_vm_group_bin_8156 (RW)
0x11e: frame_vm_group_bin_1002 (RW)
0x11f: frame_vm_group_bin_17193 (RW)
0x120: frame_vm_group_bin_9986 (RW)
0x121: frame_vm_group_bin_2828 (RW)
0x122: frame_vm_group_bin_18902 (RW)
0x123: frame_vm_group_bin_11767 (RW)
0x124: frame_vm_group_bin_4633 (RW)
0x125: frame_vm_group_bin_20754 (RW)
0x126: frame_vm_group_bin_13555 (RW)
0x127: frame_vm_group_bin_6369 (RW)
0x128: frame_vm_group_bin_22562 (RW)
0x129: frame_vm_group_bin_15380 (RW)
0x12: frame_vm_group_bin_11143 (RW)
0x12a: frame_vm_group_bin_8189 (RW)
0x12b: frame_vm_group_bin_2373 (RW)
0x12c: frame_vm_group_bin_17226 (RW)
0x12d: frame_vm_group_bin_10019 (RW)
0x12e: frame_vm_group_bin_2860 (RW)
0x12f: frame_vm_group_bin_18935 (RW)
0x130: frame_vm_group_bin_11792 (RW)
0x131: frame_vm_group_bin_4666 (RW)
0x132: frame_vm_group_bin_20787 (RW)
0x133: frame_vm_group_bin_13588 (RW)
0x134: frame_vm_group_bin_6399 (RW)
0x135: frame_vm_group_bin_22595 (RW)
0x136: frame_vm_group_bin_15413 (RW)
0x137: frame_vm_group_bin_8222 (RW)
0x138: frame_vm_group_bin_1049 (RW)
0x139: frame_vm_group_bin_17258 (RW)
0x13: frame_vm_group_bin_3958 (RW)
0x13a: frame_vm_group_bin_10053 (RW)
0x13b: frame_vm_group_bin_2896 (RW)
0x13c: frame_vm_group_bin_18967 (RW)
0x13d: frame_vm_group_bin_11825 (RW)
0x13e: frame_vm_group_bin_4698 (RW)
0x13f: frame_vm_group_bin_20820 (RW)
0x140: frame_vm_group_bin_13622 (RW)
0x141: frame_vm_group_bin_6432 (RW)
0x142: frame_vm_group_bin_22629 (RW)
0x143: frame_vm_group_bin_15447 (RW)
0x144: frame_vm_group_bin_8256 (RW)
0x145: frame_vm_group_bin_1073 (RW)
0x146: frame_vm_group_bin_17292 (RW)
0x147: frame_vm_group_bin_10086 (RW)
0x148: frame_vm_group_bin_2929 (RW)
0x149: frame_vm_group_bin_18999 (RW)
0x14: frame_vm_group_bin_20055 (RW)
0x14a: frame_vm_group_bin_11855 (RW)
0x14b: frame_vm_group_bin_4730 (RW)
0x14c: frame_vm_group_bin_1649 (RW)
0x14d: frame_vm_group_bin_13654 (RW)
0x14e: frame_vm_group_bin_6465 (RW)
0x14f: frame_vm_group_bin_22662 (RW)
0x150: frame_vm_group_bin_15480 (RW)
0x151: frame_vm_group_bin_8288 (RW)
0x152: frame_vm_group_bin_1100 (RW)
0x153: frame_vm_group_bin_17325 (RW)
0x154: frame_vm_group_bin_10119 (RW)
0x155: frame_vm_group_bin_2962 (RW)
0x156: frame_vm_group_bin_19032 (RW)
0x157: frame_vm_group_bin_11883 (RW)
0x158: frame_vm_group_bin_4763 (RW)
0x159: frame_vm_group_bin_20874 (RW)
0x15: frame_vm_group_bin_12855 (RW)
0x15a: frame_vm_group_bin_13688 (RW)
0x15b: frame_vm_group_bin_6499 (RW)
0x15c: frame_vm_group_bin_22696 (RW)
0x15d: frame_vm_group_bin_15513 (RW)
0x15e: frame_vm_group_bin_8322 (RW)
0x15f: frame_vm_group_bin_1133 (RW)
0x160: frame_vm_group_bin_17358 (RW)
0x161: frame_vm_group_bin_10155 (RW)
0x162: frame_vm_group_bin_2996 (RW)
0x163: frame_vm_group_bin_19066 (RW)
0x164: frame_vm_group_bin_11907 (RW)
0x165: frame_vm_group_bin_4797 (RW)
0x166: frame_vm_group_bin_20902 (RW)
0x167: frame_vm_group_bin_13720 (RW)
0x168: frame_vm_group_bin_6532 (RW)
0x169: frame_vm_group_bin_22729 (RW)
0x16: frame_vm_group_bin_5776 (RW)
0x16a: frame_vm_group_bin_15545 (RW)
0x16b: frame_vm_group_bin_8355 (RW)
0x16c: frame_vm_group_bin_1166 (RW)
0x16d: frame_vm_group_bin_9390 (RW)
0x16e: frame_vm_group_bin_10188 (RW)
0x16f: frame_vm_group_bin_3029 (RW)
0x170: frame_vm_group_bin_19099 (RW)
0x171: frame_vm_group_bin_11937 (RW)
0x172: frame_vm_group_bin_4829 (RW)
0x173: frame_vm_group_bin_20930 (RW)
0x174: frame_vm_group_bin_13753 (RW)
0x175: frame_vm_group_bin_6565 (RW)
0x176: frame_vm_group_bin_22761 (RW)
0x177: frame_vm_group_bin_15578 (RW)
0x178: frame_vm_group_bin_8388 (RW)
0x179: frame_vm_group_bin_1199 (RW)
0x17: frame_vm_group_bin_21892 (RW)
0x17a: frame_vm_group_bin_17417 (RW)
0x17b: frame_vm_group_bin_10222 (RW)
0x17c: frame_vm_group_bin_3063 (RW)
0x17d: frame_vm_group_bin_19131 (RW)
0x17e: frame_vm_group_bin_11968 (RW)
0x17f: frame_vm_group_bin_4863 (RW)
0x180: frame_vm_group_bin_20958 (RW)
0x181: frame_vm_group_bin_13788 (RW)
0x182: frame_vm_group_bin_6599 (RW)
0x183: frame_vm_group_bin_22795 (RW)
0x184: frame_vm_group_bin_15612 (RW)
0x185: frame_vm_group_bin_8422 (RW)
0x186: frame_vm_group_bin_1233 (RW)
0x187: frame_vm_group_bin_17441 (RW)
0x188: frame_vm_group_bin_10255 (RW)
0x189: frame_vm_group_bin_3096 (RW)
0x18: frame_vm_group_bin_14717 (RW)
0x18a: frame_vm_group_bin_19164 (RW)
0x18b: frame_vm_group_bin_12000 (RW)
0x18c: frame_vm_group_bin_4896 (RW)
0x18d: frame_vm_group_bin_20989 (RW)
0x18e: frame_vm_group_bin_13820 (RW)
0x18f: frame_vm_group_bin_6632 (RW)
0x190: frame_vm_group_bin_22828 (RW)
0x191: frame_vm_group_bin_15645 (RW)
0x192: frame_vm_group_bin_8455 (RW)
0x193: frame_vm_group_bin_1265 (RW)
0x194: frame_vm_group_bin_17463 (RW)
0x195: frame_vm_group_bin_10288 (RW)
0x196: frame_vm_group_bin_3128 (RW)
0x197: frame_vm_group_bin_19197 (RW)
0x198: frame_vm_group_bin_12030 (RW)
0x199: frame_vm_group_bin_4928 (RW)
0x19: frame_vm_group_bin_7503 (RW)
0x19a: frame_vm_group_bin_21023 (RW)
0x19b: frame_vm_group_bin_13850 (RW)
0x19c: frame_vm_group_bin_6666 (RW)
0x19d: frame_vm_group_bin_22862 (RW)
0x19e: frame_vm_group_bin_15679 (RW)
0x19f: frame_vm_group_bin_8489 (RW)
0x1: frame_vm_group_bin_16466 (RW)
0x1a0: frame_vm_group_bin_1297 (RW)
0x1a1: frame_vm_group_bin_17484 (RW)
0x1a2: frame_vm_group_bin_10322 (RW)
0x1a3: frame_vm_group_bin_3162 (RW)
0x1a4: frame_vm_group_bin_19231 (RW)
0x1a5: frame_vm_group_bin_12059 (RW)
0x1a6: frame_vm_group_bin_4960 (RW)
0x1a7: frame_vm_group_bin_21057 (RW)
0x1a8: frame_vm_group_bin_13879 (RW)
0x1a9: frame_vm_group_bin_6699 (RW)
0x1a: frame_vm_group_bin_0349 (RW)
0x1aa: frame_vm_group_bin_22895 (RW)
0x1ab: frame_vm_group_bin_15712 (RW)
0x1ac: frame_vm_group_bin_8521 (RW)
0x1ad: frame_vm_group_bin_1329 (RW)
0x1ae: frame_vm_group_bin_17508 (RW)
0x1af: frame_vm_group_bin_10355 (RW)
0x1b0: frame_vm_group_bin_3195 (RW)
0x1b1: frame_vm_group_bin_19264 (RW)
0x1b2: frame_vm_group_bin_12091 (RW)
0x1b3: frame_vm_group_bin_4992 (RW)
0x1b4: frame_vm_group_bin_21090 (RW)
0x1b5: frame_vm_group_bin_13912 (RW)
0x1b6: frame_vm_group_bin_6731 (RW)
0x1b7: frame_vm_group_bin_22928 (RW)
0x1b8: frame_vm_group_bin_15745 (RW)
0x1b9: frame_vm_group_bin_8553 (RW)
0x1b: frame_vm_group_bin_16533 (RW)
0x1ba: frame_vm_group_bin_1365 (RW)
0x1bb: frame_vm_group_bin_17537 (RW)
0x1bc: frame_vm_group_bin_10388 (RW)
0x1bd: frame_vm_group_bin_3229 (RW)
0x1be: frame_vm_group_bin_19298 (RW)
0x1bf: frame_vm_group_bin_12124 (RW)
0x1c0: frame_vm_group_bin_5026 (RW)
0x1c1: frame_vm_group_bin_21124 (RW)
0x1c2: frame_vm_group_bin_13946 (RW)
0x1c3: frame_vm_group_bin_6764 (RW)
0x1c4: frame_vm_group_bin_22961 (RW)
0x1c5: frame_vm_group_bin_15779 (RW)
0x1c6: frame_vm_group_bin_8586 (RW)
0x1c7: frame_vm_group_bin_1397 (RW)
0x1c8: frame_vm_group_bin_17558 (RW)
0x1c9: frame_vm_group_bin_10413 (RW)
0x1c: frame_vm_group_bin_9321 (RW)
0x1ca: frame_vm_group_bin_3261 (RW)
0x1cb: frame_vm_group_bin_19331 (RW)
0x1cc: frame_vm_group_bin_12157 (RW)
0x1cd: frame_vm_group_bin_5059 (RW)
0x1ce: frame_vm_group_bin_21156 (RW)
0x1cf: frame_vm_group_bin_13979 (RW)
0x1d0: frame_vm_group_bin_6797 (RW)
0x1d1: frame_vm_group_bin_22994 (RW)
0x1d2: frame_vm_group_bin_15811 (RW)
0x1d3: frame_vm_group_bin_8618 (RW)
0x1d4: frame_vm_group_bin_1430 (RW)
0x1d5: frame_vm_group_bin_17581 (RW)
0x1d6: frame_vm_group_bin_10441 (RW)
0x1d7: frame_vm_group_bin_3294 (RW)
0x1d8: frame_vm_group_bin_19364 (RW)
0x1d9: frame_vm_group_bin_12186 (RW)
0x1d: frame_vm_group_bin_2171 (RW)
0x1da: frame_vm_group_bin_5094 (RW)
0x1db: frame_vm_group_bin_21190 (RW)
0x1dc: frame_vm_group_bin_14013 (RW)
0x1dd: frame_vm_group_bin_6828 (RW)
0x1de: frame_vm_group_bin_23027 (RW)
0x1df: frame_vm_group_bin_15844 (RW)
0x1e0: frame_vm_group_bin_8652 (RW)
0x1e1: frame_vm_group_bin_1464 (RW)
0x1e2: frame_vm_group_bin_17606 (RW)
0x1e3: frame_vm_group_bin_10475 (RW)
0x1e4: frame_vm_group_bin_3328 (RW)
0x1e5: frame_vm_group_bin_19398 (RW)
0x1e6: frame_vm_group_bin_12217 (RW)
0x1e7: frame_vm_group_bin_5127 (RW)
0x1e8: frame_vm_group_bin_21223 (RW)
0x1e9: frame_vm_group_bin_14046 (RW)
0x1e: frame_vm_group_bin_18265 (RW)
0x1ea: frame_vm_group_bin_6855 (RW)
0x1eb: frame_vm_group_bin_23060 (RW)
0x1ec: frame_vm_group_bin_15877 (RW)
0x1ed: frame_vm_group_bin_8686 (RW)
0x1ee: frame_vm_group_bin_1497 (RW)
0x1ef: frame_vm_group_bin_17637 (RW)
0x1f0: frame_vm_group_bin_10508 (RW)
0x1f1: frame_vm_group_bin_3361 (RW)
0x1f2: frame_vm_group_bin_19430 (RW)
0x1f3: frame_vm_group_bin_12249 (RW)
0x1f4: frame_vm_group_bin_5160 (RW)
0x1f5: frame_vm_group_bin_21256 (RW)
0x1f6: frame_vm_group_bin_14079 (RW)
0x1f7: frame_vm_group_bin_6880 (RW)
0x1f8: frame_vm_group_bin_23093 (RW)
0x1f9: frame_vm_group_bin_15910 (RW)
0x1f: frame_vm_group_bin_11177 (RW)
0x1fa: frame_vm_group_bin_8720 (RW)
0x1fb: frame_vm_group_bin_1531 (RW)
0x1fc: frame_vm_group_bin_17671 (RW)
0x1fd: frame_vm_group_bin_10541 (RW)
0x1fe: frame_vm_group_bin_3392 (RW)
0x1ff: frame_vm_group_bin_19461 (RW)
0x20: frame_vm_group_bin_3992 (RW)
0x21: frame_vm_group_bin_20089 (RW)
0x22: frame_vm_group_bin_12889 (RW)
0x23: frame_vm_group_bin_7996 (RW)
0x24: frame_vm_group_bin_21925 (RW)
0x25: frame_vm_group_bin_14750 (RW)
0x26: frame_vm_group_bin_7535 (RW)
0x27: frame_vm_group_bin_0381 (RW)
0x28: frame_vm_group_bin_16565 (RW)
0x29: frame_vm_group_bin_9354 (RW)
0x2: frame_vm_group_bin_9264 (RW)
0x2a: frame_vm_group_bin_21284 (RW)
0x2b: frame_vm_group_bin_18298 (RW)
0x2c: frame_vm_group_bin_11210 (RW)
0x2d: frame_vm_group_bin_4025 (RW)
0x2e: frame_vm_group_bin_20121 (RW)
0x2f: frame_vm_group_bin_12922 (RW)
0x30: frame_vm_group_bin_5820 (RW)
0x31: frame_vm_group_bin_21958 (RW)
0x32: frame_vm_group_bin_14782 (RW)
0x33: frame_vm_group_bin_7567 (RW)
0x34: frame_vm_group_bin_0409 (RW)
0x35: frame_vm_group_bin_16597 (RW)
0x36: frame_vm_group_bin_9387 (RW)
0x37: frame_vm_group_bin_2230 (RW)
0x38: frame_vm_group_bin_18331 (RW)
0x39: frame_vm_group_bin_11243 (RW)
0x3: frame_vm_group_bin_2103 (RW)
0x3a: frame_vm_group_bin_4059 (RW)
0x3b: frame_vm_group_bin_20155 (RW)
0x3c: frame_vm_group_bin_12955 (RW)
0x3d: frame_vm_group_bin_5846 (RW)
0x3e: frame_vm_group_bin_21992 (RW)
0x3f: frame_vm_group_bin_14816 (RW)
0x40: frame_vm_group_bin_7601 (RW)
0x41: frame_vm_group_bin_0441 (RW)
0x42: frame_vm_group_bin_16631 (RW)
0x43: frame_vm_group_bin_9422 (RW)
0x44: frame_vm_group_bin_2262 (RW)
0x45: frame_vm_group_bin_18365 (RW)
0x46: frame_vm_group_bin_11277 (RW)
0x47: frame_vm_group_bin_4092 (RW)
0x48: frame_vm_group_bin_20186 (RW)
0x49: frame_vm_group_bin_12988 (RW)
0x4: frame_vm_group_bin_18198 (RW)
0x4a: frame_vm_group_bin_5871 (RW)
0x4b: frame_vm_group_bin_7927 (RW)
0x4c: frame_vm_group_bin_14849 (RW)
0x4d: frame_vm_group_bin_7634 (RW)
0x4e: frame_vm_group_bin_0474 (RW)
0x4f: frame_vm_group_bin_16664 (RW)
0x50: frame_vm_group_bin_9455 (RW)
0x51: frame_vm_group_bin_2295 (RW)
0x52: frame_vm_group_bin_18397 (RW)
0x53: frame_vm_group_bin_11310 (RW)
0x54: frame_vm_group_bin_4124 (RW)
0x55: frame_vm_group_bin_20219 (RW)
0x56: frame_vm_group_bin_13023 (RW)
0x57: frame_vm_group_bin_5896 (RW)
0x58: frame_vm_group_bin_22044 (RW)
0x59: frame_vm_group_bin_14882 (RW)
0x5: frame_vm_group_bin_11111 (RW)
0x5a: frame_vm_group_bin_7668 (RW)
0x5b: frame_vm_group_bin_0507 (RW)
0x5c: frame_vm_group_bin_16697 (RW)
0x5d: frame_vm_group_bin_9489 (RW)
0x5e: frame_vm_group_bin_2329 (RW)
0x5f: frame_vm_group_bin_18430 (RW)
0x60: frame_vm_group_bin_11342 (RW)
0x61: frame_vm_group_bin_4157 (RW)
0x62: frame_vm_group_bin_20253 (RW)
0x63: frame_vm_group_bin_13057 (RW)
0x64: frame_vm_group_bin_5924 (RW)
0x65: frame_vm_group_bin_22068 (RW)
0x66: frame_vm_group_bin_14916 (RW)
0x67: frame_vm_group_bin_7701 (RW)
0x68: frame_vm_group_bin_0539 (RW)
0x69: frame_vm_group_bin_16731 (RW)
0x6: frame_vm_group_bin_3926 (RW)
0x6a: frame_vm_group_bin_9522 (RW)
0x6b: frame_vm_group_bin_2362 (RW)
0x6c: frame_vm_group_bin_18462 (RW)
0x6d: frame_vm_group_bin_11375 (RW)
0x6e: frame_vm_group_bin_4190 (RW)
0x6f: frame_vm_group_bin_20285 (RW)
0x70: frame_vm_group_bin_13090 (RW)
0x71: frame_vm_group_bin_5946 (RW)
0x72: frame_vm_group_bin_22098 (RW)
0x73: frame_vm_group_bin_14949 (RW)
0x74: frame_vm_group_bin_7733 (RW)
0x75: frame_vm_group_bin_0570 (RW)
0x76: frame_vm_group_bin_16764 (RW)
0x77: frame_vm_group_bin_9555 (RW)
0x78: frame_vm_group_bin_2395 (RW)
0x79: frame_vm_group_bin_18489 (RW)
0x7: frame_vm_group_bin_20022 (RW)
0x7a: frame_vm_group_bin_11408 (RW)
0x7b: frame_vm_group_bin_4223 (RW)
0x7c: frame_vm_group_bin_20321 (RW)
0x7d: frame_vm_group_bin_13124 (RW)
0x7e: frame_vm_group_bin_5971 (RW)
0x7f: frame_vm_group_bin_22132 (RW)
0x80: frame_vm_group_bin_14983 (RW)
0x81: frame_vm_group_bin_7767 (RW)
0x82: frame_vm_group_bin_0603 (RW)
0x83: frame_vm_group_bin_16798 (RW)
0x84: frame_vm_group_bin_9589 (RW)
0x85: frame_vm_group_bin_2428 (RW)
0x86: frame_vm_group_bin_18517 (RW)
0x87: frame_vm_group_bin_11440 (RW)
0x88: frame_vm_group_bin_4256 (RW)
0x89: frame_vm_group_bin_20354 (RW)
0x8: frame_vm_group_bin_12822 (RW)
0x8a: frame_vm_group_bin_13157 (RW)
0x8b: frame_vm_group_bin_6002 (RW)
0x8c: frame_vm_group_bin_22165 (RW)
0x8d: frame_vm_group_bin_15016 (RW)
0x8e: frame_vm_group_bin_7800 (RW)
0x8f: frame_vm_group_bin_0634 (RW)
0x90: frame_vm_group_bin_16831 (RW)
0x91: frame_vm_group_bin_9622 (RW)
0x92: frame_vm_group_bin_2461 (RW)
0x93: frame_vm_group_bin_18541 (RW)
0x94: frame_vm_group_bin_11473 (RW)
0x95: frame_vm_group_bin_4289 (RW)
0x96: frame_vm_group_bin_20387 (RW)
0x97: frame_vm_group_bin_13190 (RW)
0x98: frame_vm_group_bin_6033 (RW)
0x99: frame_vm_group_bin_22198 (RW)
0x9: frame_vm_group_bin_22010 (RW)
0x9a: frame_vm_group_bin_15045 (RW)
0x9b: frame_vm_group_bin_7833 (RW)
0x9c: frame_vm_group_bin_0669 (RW)
0x9d: frame_vm_group_bin_19505 (RW)
0x9e: frame_vm_group_bin_9656 (RW)
0x9f: frame_vm_group_bin_2494 (RW)
0xa0: frame_vm_group_bin_18571 (RW)
0xa1: frame_vm_group_bin_11507 (RW)
0xa2: frame_vm_group_bin_4323 (RW)
0xa3: frame_vm_group_bin_20421 (RW)
0xa4: frame_vm_group_bin_13224 (RW)
0xa5: frame_vm_group_bin_6059 (RW)
0xa6: frame_vm_group_bin_22232 (RW)
0xa7: frame_vm_group_bin_15069 (RW)
0xa8: frame_vm_group_bin_7866 (RW)
0xa9: frame_vm_group_bin_0702 (RW)
0xa: frame_vm_group_bin_21859 (RW)
0xaa: frame_vm_group_bin_16896 (RW)
0xab: frame_vm_group_bin_9688 (RW)
0xac: frame_vm_group_bin_2527 (RW)
0xad: frame_vm_group_bin_18604 (RW)
0xae: frame_vm_group_bin_11540 (RW)
0xaf: frame_vm_group_bin_4358 (RW)
0xb0: frame_vm_group_bin_20454 (RW)
0xb1: frame_vm_group_bin_13257 (RW)
0xb2: frame_vm_group_bin_6085 (RW)
0xb3: frame_vm_group_bin_22265 (RW)
0xb4: frame_vm_group_bin_15093 (RW)
0xb5: frame_vm_group_bin_7899 (RW)
0xb6: frame_vm_group_bin_0735 (RW)
0xb7: frame_vm_group_bin_16929 (RW)
0xb8: frame_vm_group_bin_9721 (RW)
0xb9: frame_vm_group_bin_2560 (RW)
0xb: frame_vm_group_bin_14684 (RW)
0xba: frame_vm_group_bin_1224 (RW)
0xbb: frame_vm_group_bin_11571 (RW)
0xbc: frame_vm_group_bin_4392 (RW)
0xbd: frame_vm_group_bin_20488 (RW)
0xbe: frame_vm_group_bin_13291 (RW)
0xbf: frame_vm_group_bin_6116 (RW)
0xc0: frame_vm_group_bin_22298 (RW)
0xc1: frame_vm_group_bin_15123 (RW)
0xc2: frame_vm_group_bin_7934 (RW)
0xc3: frame_vm_group_bin_0769 (RW)
0xc4: frame_vm_group_bin_16963 (RW)
0xc5: frame_vm_group_bin_9755 (RW)
0xc6: frame_vm_group_bin_2594 (RW)
0xc7: frame_vm_group_bin_18670 (RW)
0xc8: frame_vm_group_bin_11596 (RW)
0xc9: frame_vm_group_bin_4425 (RW)
0xc: frame_vm_group_bin_7470 (RW)
0xca: frame_vm_group_bin_20521 (RW)
0xcb: frame_vm_group_bin_13323 (RW)
0xcc: frame_vm_group_bin_6148 (RW)
0xcd: frame_vm_group_bin_22331 (RW)
0xce: frame_vm_group_bin_15146 (RW)
0xcf: frame_vm_group_bin_7967 (RW)
0xd0: frame_vm_group_bin_0802 (RW)
0xd1: frame_vm_group_bin_16996 (RW)
0xd2: frame_vm_group_bin_9788 (RW)
0xd3: frame_vm_group_bin_2627 (RW)
0xd4: frame_vm_group_bin_18702 (RW)
0xd5: frame_vm_group_bin_11621 (RW)
0xd6: frame_vm_group_bin_4458 (RW)
0xd7: frame_vm_group_bin_20554 (RW)
0xd8: frame_vm_group_bin_13356 (RW)
0xd9: frame_vm_group_bin_6181 (RW)
0xd: frame_vm_group_bin_0317 (RW)
0xda: frame_vm_group_bin_22364 (RW)
0xdb: frame_vm_group_bin_15180 (RW)
0xdc: frame_vm_group_bin_7999 (RW)
0xdd: frame_vm_group_bin_0835 (RW)
0xde: frame_vm_group_bin_17030 (RW)
0xdf: frame_vm_group_bin_9822 (RW)
0xe0: frame_vm_group_bin_2661 (RW)
0xe1: frame_vm_group_bin_18734 (RW)
0xe2: frame_vm_group_bin_11645 (RW)
0xe3: frame_vm_group_bin_4492 (RW)
0xe4: frame_vm_group_bin_20588 (RW)
0xe5: frame_vm_group_bin_13388 (RW)
0xe6: frame_vm_group_bin_6210 (RW)
0xe7: frame_vm_group_bin_22397 (RW)
0xe8: frame_vm_group_bin_15213 (RW)
0xe9: frame_vm_group_bin_8027 (RW)
0xe: frame_vm_group_bin_16499 (RW)
0xea: frame_vm_group_bin_0868 (RW)
0xeb: frame_vm_group_bin_17063 (RW)
0xec: frame_vm_group_bin_9855 (RW)
0xed: frame_vm_group_bin_2694 (RW)
0xee: frame_vm_group_bin_18767 (RW)
0xef: frame_vm_group_bin_11666 (RW)
0xf0: frame_vm_group_bin_4525 (RW)
0xf1: frame_vm_group_bin_20621 (RW)
0xf2: frame_vm_group_bin_13421 (RW)
0xf3: frame_vm_group_bin_6238 (RW)
0xf4: frame_vm_group_bin_22429 (RW)
0xf5: frame_vm_group_bin_15247 (RW)
0xf6: frame_vm_group_bin_8057 (RW)
0xf7: frame_vm_group_bin_0901 (RW)
0xf8: frame_vm_group_bin_17096 (RW)
0xf9: frame_vm_group_bin_4176 (RW)
0xf: frame_vm_group_bin_9290 (RW)
0xfa: frame_vm_group_bin_2728 (RW)
0xfb: frame_vm_group_bin_18801 (RW)
0xfc: frame_vm_group_bin_11693 (RW)
0xfd: frame_vm_group_bin_4558 (RW)
0xfe: frame_vm_group_bin_20654 (RW)
0xff: frame_vm_group_bin_13455 (RW)
}
pt_vm_group_bin_0380 {
0x0: frame_vm_group_bin_2125 (RW)
0x100: frame_vm_group_bin_8110 (RW)
0x101: frame_vm_group_bin_0956 (RW)
0x102: frame_vm_group_bin_17150 (RW)
0x103: frame_vm_group_bin_9940 (RW)
0x104: frame_vm_group_bin_2782 (RW)
0x105: frame_vm_group_bin_18856 (RW)
0x106: frame_vm_group_bin_20461 (RW)
0x107: frame_vm_group_bin_4599 (RW)
0x108: frame_vm_group_bin_20708 (RW)
0x109: frame_vm_group_bin_13509 (RW)
0x10: frame_vm_group_bin_3979 (RW)
0x10a: frame_vm_group_bin_6323 (RW)
0x10b: frame_vm_group_bin_22517 (RW)
0x10c: frame_vm_group_bin_15334 (RW)
0x10d: frame_vm_group_bin_8143 (RW)
0x10e: frame_vm_group_bin_0989 (RW)
0x10f: frame_vm_group_bin_17182 (RW)
0x110: frame_vm_group_bin_9973 (RW)
0x111: frame_vm_group_bin_2815 (RW)
0x112: frame_vm_group_bin_18889 (RW)
0x113: frame_vm_group_bin_11756 (RW)
0x114: frame_vm_group_bin_4623 (RW)
0x115: frame_vm_group_bin_20741 (RW)
0x116: frame_vm_group_bin_13542 (RW)
0x117: frame_vm_group_bin_6356 (RW)
0x118: frame_vm_group_bin_22549 (RW)
0x119: frame_vm_group_bin_15367 (RW)
0x11: frame_vm_group_bin_20076 (RW)
0x11a: frame_vm_group_bin_8177 (RW)
0x11b: frame_vm_group_bin_1020 (RW)
0x11c: frame_vm_group_bin_17214 (RW)
0x11d: frame_vm_group_bin_10007 (RW)
0x11e: frame_vm_group_bin_2849 (RW)
0x11f: frame_vm_group_bin_18923 (RW)
0x120: frame_vm_group_bin_6452 (RW)
0x121: frame_vm_group_bin_4654 (RW)
0x122: frame_vm_group_bin_20775 (RW)
0x123: frame_vm_group_bin_13576 (RW)
0x124: frame_vm_group_bin_6387 (RW)
0x125: frame_vm_group_bin_22583 (RW)
0x126: frame_vm_group_bin_15401 (RW)
0x127: frame_vm_group_bin_8210 (RW)
0x128: frame_vm_group_bin_1043 (RW)
0x129: frame_vm_group_bin_17246 (RW)
0x12: frame_vm_group_bin_12876 (RW)
0x12a: frame_vm_group_bin_10040 (RW)
0x12b: frame_vm_group_bin_2883 (RW)
0x12c: frame_vm_group_bin_18955 (RW)
0x12d: frame_vm_group_bin_11812 (RW)
0x12e: frame_vm_group_bin_4686 (RW)
0x12f: frame_vm_group_bin_20808 (RW)
0x130: frame_vm_group_bin_13609 (RW)
0x131: frame_vm_group_bin_6419 (RW)
0x132: frame_vm_group_bin_22616 (RW)
0x133: frame_vm_group_bin_15434 (RW)
0x134: frame_vm_group_bin_8243 (RW)
0x135: frame_vm_group_bin_1064 (RW)
0x136: frame_vm_group_bin_17279 (RW)
0x137: frame_vm_group_bin_10073 (RW)
0x138: frame_vm_group_bin_2916 (RW)
0x139: frame_vm_group_bin_18986 (RW)
0x13: frame_vm_group_bin_5792 (RW)
0x13a: frame_vm_group_bin_15838 (RW)
0x13b: frame_vm_group_bin_4719 (RW)
0x13c: frame_vm_group_bin_20841 (RW)
0x13d: frame_vm_group_bin_13642 (RW)
0x13e: frame_vm_group_bin_6454 (RW)
0x13f: frame_vm_group_bin_22650 (RW)
0x140: frame_vm_group_bin_15468 (RW)
0x141: frame_vm_group_bin_8276 (RW)
0x142: frame_vm_group_bin_1092 (RW)
0x143: frame_vm_group_bin_17313 (RW)
0x144: frame_vm_group_bin_10107 (RW)
0x145: frame_vm_group_bin_2950 (RW)
0x146: frame_vm_group_bin_19020 (RW)
0x147: frame_vm_group_bin_11873 (RW)
0x148: frame_vm_group_bin_4751 (RW)
0x149: frame_vm_group_bin_20866 (RW)
0x14: frame_vm_group_bin_21913 (RW)
0x14a: frame_vm_group_bin_13675 (RW)
0x14b: frame_vm_group_bin_6486 (RW)
0x14c: frame_vm_group_bin_22683 (RW)
0x14d: frame_vm_group_bin_15501 (RW)
0x14e: frame_vm_group_bin_8309 (RW)
0x14f: frame_vm_group_bin_1120 (RW)
0x150: frame_vm_group_bin_17346 (RW)
0x151: frame_vm_group_bin_10140 (RW)
0x152: frame_vm_group_bin_2983 (RW)
0x153: frame_vm_group_bin_19053 (RW)
0x154: frame_vm_group_bin_1835 (RW)
0x155: frame_vm_group_bin_4784 (RW)
0x156: frame_vm_group_bin_20892 (RW)
0x157: frame_vm_group_bin_13708 (RW)
0x158: frame_vm_group_bin_6519 (RW)
0x159: frame_vm_group_bin_22716 (RW)
0x15: frame_vm_group_bin_14737 (RW)
0x15a: frame_vm_group_bin_15534 (RW)
0x15b: frame_vm_group_bin_8343 (RW)
0x15c: frame_vm_group_bin_1154 (RW)
0x15d: frame_vm_group_bin_17379 (RW)
0x15e: frame_vm_group_bin_10176 (RW)
0x15f: frame_vm_group_bin_3017 (RW)
0x160: frame_vm_group_bin_19087 (RW)
0x161: frame_vm_group_bin_11925 (RW)
0x162: frame_vm_group_bin_4817 (RW)
0x163: frame_vm_group_bin_20921 (RW)
0x164: frame_vm_group_bin_13741 (RW)
0x165: frame_vm_group_bin_6553 (RW)
0x166: frame_vm_group_bin_22749 (RW)
0x167: frame_vm_group_bin_15566 (RW)
0x168: frame_vm_group_bin_8376 (RW)
0x169: frame_vm_group_bin_1187 (RW)
0x16: frame_vm_group_bin_7523 (RW)
0x16a: frame_vm_group_bin_17407 (RW)
0x16b: frame_vm_group_bin_10209 (RW)
0x16c: frame_vm_group_bin_3050 (RW)
0x16d: frame_vm_group_bin_19119 (RW)
0x16e: frame_vm_group_bin_11955 (RW)
0x16f: frame_vm_group_bin_4850 (RW)
0x170: frame_vm_group_bin_20948 (RW)
0x171: frame_vm_group_bin_13775 (RW)
0x172: frame_vm_group_bin_6586 (RW)
0x173: frame_vm_group_bin_22782 (RW)
0x174: frame_vm_group_bin_15599 (RW)
0x175: frame_vm_group_bin_8409 (RW)
0x176: frame_vm_group_bin_1220 (RW)
0x177: frame_vm_group_bin_17431 (RW)
0x178: frame_vm_group_bin_10242 (RW)
0x179: frame_vm_group_bin_3083 (RW)
0x17: frame_vm_group_bin_0369 (RW)
0x17a: frame_vm_group_bin_19152 (RW)
0x17b: frame_vm_group_bin_11989 (RW)
0x17c: frame_vm_group_bin_4884 (RW)
0x17d: frame_vm_group_bin_20977 (RW)
0x17e: frame_vm_group_bin_13809 (RW)
0x17f: frame_vm_group_bin_6620 (RW)
0x180: frame_vm_group_bin_22816 (RW)
0x181: frame_vm_group_bin_15633 (RW)
0x182: frame_vm_group_bin_8443 (RW)
0x183: frame_vm_group_bin_1253 (RW)
0x184: frame_vm_group_bin_2965 (RW)
0x185: frame_vm_group_bin_10276 (RW)
0x186: frame_vm_group_bin_3116 (RW)
0x187: frame_vm_group_bin_19185 (RW)
0x188: frame_vm_group_bin_12020 (RW)
0x189: frame_vm_group_bin_4917 (RW)
0x18: frame_vm_group_bin_12096 (RW)
0x18a: frame_vm_group_bin_21010 (RW)
0x18b: frame_vm_group_bin_13838 (RW)
0x18c: frame_vm_group_bin_6653 (RW)
0x18d: frame_vm_group_bin_22849 (RW)
0x18e: frame_vm_group_bin_15666 (RW)
0x18f: frame_vm_group_bin_8476 (RW)
0x190: frame_vm_group_bin_1284 (RW)
0x191: frame_vm_group_bin_7571 (RW)
0x192: frame_vm_group_bin_10309 (RW)
0x193: frame_vm_group_bin_3149 (RW)
0x194: frame_vm_group_bin_19218 (RW)
0x195: frame_vm_group_bin_1859 (RW)
0x196: frame_vm_group_bin_4948 (RW)
0x197: frame_vm_group_bin_21043 (RW)
0x198: frame_vm_group_bin_13867 (RW)
0x199: frame_vm_group_bin_6686 (RW)
0x19: frame_vm_group_bin_9341 (RW)
0x19a: frame_vm_group_bin_22883 (RW)
0x19b: frame_vm_group_bin_15700 (RW)
0x19c: frame_vm_group_bin_8510 (RW)
0x19d: frame_vm_group_bin_1317 (RW)
0x19e: frame_vm_group_bin_12230 (RW)
0x19f: frame_vm_group_bin_10343 (RW)
0x1: frame_vm_group_bin_18219 (RW)
0x1a0: frame_vm_group_bin_3183 (RW)
0x1a1: frame_vm_group_bin_19252 (RW)
0x1a2: frame_vm_group_bin_12079 (RW)
0x1a3: frame_vm_group_bin_4980 (RW)
0x1a4: frame_vm_group_bin_21078 (RW)
0x1a5: frame_vm_group_bin_13900 (RW)
0x1a6: frame_vm_group_bin_6719 (RW)
0x1a7: frame_vm_group_bin_22916 (RW)
0x1a8: frame_vm_group_bin_15733 (RW)
0x1a9: frame_vm_group_bin_8542 (RW)
0x1a: frame_vm_group_bin_2191 (RW)
0x1aa: frame_vm_group_bin_1350 (RW)
0x1ab: frame_vm_group_bin_16979 (RW)
0x1ac: frame_vm_group_bin_10376 (RW)
0x1ad: frame_vm_group_bin_3216 (RW)
0x1ae: frame_vm_group_bin_19285 (RW)
0x1af: frame_vm_group_bin_11244 (RW)
0x1b0: frame_vm_group_bin_5013 (RW)
0x1b1: frame_vm_group_bin_21111 (RW)
0x1b2: frame_vm_group_bin_13933 (RW)
0x1b3: frame_vm_group_bin_6752 (RW)
0x1b4: frame_vm_group_bin_22949 (RW)
0x1b5: frame_vm_group_bin_15766 (RW)
0x1b6: frame_vm_group_bin_8573 (RW)
0x1b7: frame_vm_group_bin_1384 (RW)
0x1b8: frame_vm_group_bin_21611 (RW)
0x1b9: frame_vm_group_bin_10403 (RW)
0x1b: frame_vm_group_bin_18286 (RW)
0x1ba: frame_vm_group_bin_3249 (RW)
0x1bb: frame_vm_group_bin_19319 (RW)
0x1bc: frame_vm_group_bin_12145 (RW)
0x1bd: frame_vm_group_bin_5047 (RW)
0x1be: frame_vm_group_bin_21144 (RW)
0x1bf: frame_vm_group_bin_13967 (RW)
0x1c0: frame_vm_group_bin_6785 (RW)
0x1c1: frame_vm_group_bin_22982 (RW)
0x1c2: frame_vm_group_bin_15799 (RW)
0x1c3: frame_vm_group_bin_8606 (RW)
0x1c4: frame_vm_group_bin_1418 (RW)
0x1c5: frame_vm_group_bin_2990 (RW)
0x1c6: frame_vm_group_bin_10432 (RW)
0x1c7: frame_vm_group_bin_3282 (RW)
0x1c8: frame_vm_group_bin_19352 (RW)
0x1c9: frame_vm_group_bin_12175 (RW)
0x1c: frame_vm_group_bin_11198 (RW)
0x1ca: frame_vm_group_bin_5081 (RW)
0x1cb: frame_vm_group_bin_21177 (RW)
0x1cc: frame_vm_group_bin_14000 (RW)
0x1cd: frame_vm_group_bin_6816 (RW)
0x1ce: frame_vm_group_bin_23014 (RW)
0x1cf: frame_vm_group_bin_15831 (RW)
0x1d0: frame_vm_group_bin_8639 (RW)
0x1d1: frame_vm_group_bin_1451 (RW)
0x1d2: frame_vm_group_bin_7595 (RW)
0x1d3: frame_vm_group_bin_10462 (RW)
0x1d4: frame_vm_group_bin_3315 (RW)
0x1d5: frame_vm_group_bin_19385 (RW)
0x1d6: frame_vm_group_bin_1882 (RW)
0x1d7: frame_vm_group_bin_5114 (RW)
0x1d8: frame_vm_group_bin_21210 (RW)
0x1d9: frame_vm_group_bin_14033 (RW)
0x1d: frame_vm_group_bin_4013 (RW)
0x1da: frame_vm_group_bin_6845 (RW)
0x1db: frame_vm_group_bin_23048 (RW)
0x1dc: frame_vm_group_bin_15865 (RW)
0x1dd: frame_vm_group_bin_8675 (RW)
0x1de: frame_vm_group_bin_1485 (RW)
0x1df: frame_vm_group_bin_17625 (RW)
0x1e0: frame_vm_group_bin_10496 (RW)
0x1e1: frame_vm_group_bin_3349 (RW)
0x1e2: frame_vm_group_bin_19418 (RW)
0x1e3: frame_vm_group_bin_12237 (RW)
0x1e4: frame_vm_group_bin_5148 (RW)
0x1e5: frame_vm_group_bin_21244 (RW)
0x1e6: frame_vm_group_bin_14067 (RW)
0x1e7: frame_vm_group_bin_6873 (RW)
0x1e8: frame_vm_group_bin_23081 (RW)
0x1e9: frame_vm_group_bin_15898 (RW)
0x1e: frame_vm_group_bin_20109 (RW)
0x1ea: frame_vm_group_bin_8707 (RW)
0x1eb: frame_vm_group_bin_1518 (RW)
0x1ec: frame_vm_group_bin_17658 (RW)
0x1ed: frame_vm_group_bin_10528 (RW)
0x1ee: frame_vm_group_bin_3380 (RW)
0x1ef: frame_vm_group_bin_19449 (RW)
0x1f0: frame_vm_group_bin_12270 (RW)
0x1f1: frame_vm_group_bin_5181 (RW)
0x1f2: frame_vm_group_bin_21277 (RW)
0x1f3: frame_vm_group_bin_14100 (RW)
0x1f4: frame_vm_group_bin_6896 (RW)
0x1f5: frame_vm_group_bin_23114 (RW)
0x1f6: frame_vm_group_bin_15931 (RW)
0x1f7: frame_vm_group_bin_8740 (RW)
0x1f8: frame_vm_group_bin_1551 (RW)
0x1f9: frame_vm_group_bin_17688 (RW)
0x1f: frame_vm_group_bin_12910 (RW)
0x1fa: frame_vm_group_bin_10562 (RW)
0x1fb: frame_vm_group_bin_3408 (RW)
0x1fc: frame_vm_group_bin_19482 (RW)
0x1fd: frame_vm_group_bin_12304 (RW)
0x1fe: frame_vm_group_bin_5215 (RW)
0x1ff: frame_vm_group_bin_21310 (RW)
0x20: frame_vm_group_bin_0643 (RW)
0x21: frame_vm_group_bin_21946 (RW)
0x22: frame_vm_group_bin_14771 (RW)
0x23: frame_vm_group_bin_7555 (RW)
0x24: frame_vm_group_bin_18191 (RW)
0x25: frame_vm_group_bin_16586 (RW)
0x26: frame_vm_group_bin_9375 (RW)
0x27: frame_vm_group_bin_2221 (RW)
0x28: frame_vm_group_bin_18319 (RW)
0x29: frame_vm_group_bin_11231 (RW)
0x2: frame_vm_group_bin_11131 (RW)
0x2a: frame_vm_group_bin_4046 (RW)
0x2b: frame_vm_group_bin_20142 (RW)
0x2c: frame_vm_group_bin_12942 (RW)
0x2d: frame_vm_group_bin_5375 (RW)
0x2e: frame_vm_group_bin_21979 (RW)
0x2f: frame_vm_group_bin_14803 (RW)
0x30: frame_vm_group_bin_7588 (RW)
0x31: frame_vm_group_bin_0428 (RW)
0x32: frame_vm_group_bin_16618 (RW)
0x33: frame_vm_group_bin_9409 (RW)
0x34: frame_vm_group_bin_2249 (RW)
0x35: frame_vm_group_bin_18352 (RW)
0x36: frame_vm_group_bin_11264 (RW)
0x37: frame_vm_group_bin_4079 (RW)
0x38: frame_vm_group_bin_20174 (RW)
0x39: frame_vm_group_bin_12975 (RW)
0x3: frame_vm_group_bin_3946 (RW)
0x3a: frame_vm_group_bin_10005 (RW)
0x3b: frame_vm_group_bin_22012 (RW)
0x3c: frame_vm_group_bin_14837 (RW)
0x3d: frame_vm_group_bin_7622 (RW)
0x3e: frame_vm_group_bin_0462 (RW)
0x3f: frame_vm_group_bin_16652 (RW)
0x40: frame_vm_group_bin_9443 (RW)
0x41: frame_vm_group_bin_2283 (RW)
0x42: frame_vm_group_bin_18386 (RW)
0x43: frame_vm_group_bin_11298 (RW)
0x44: frame_vm_group_bin_4112 (RW)
0x45: frame_vm_group_bin_20207 (RW)
0x46: frame_vm_group_bin_13011 (RW)
0x47: frame_vm_group_bin_14670 (RW)
0x48: frame_vm_group_bin_22038 (RW)
0x49: frame_vm_group_bin_14870 (RW)
0x4: frame_vm_group_bin_20043 (RW)
0x4a: frame_vm_group_bin_7655 (RW)
0x4b: frame_vm_group_bin_0494 (RW)
0x4c: frame_vm_group_bin_16685 (RW)
0x4d: frame_vm_group_bin_9476 (RW)
0x4e: frame_vm_group_bin_2316 (RW)
0x4f: frame_vm_group_bin_18417 (RW)
0x50: frame_vm_group_bin_11331 (RW)
0x51: frame_vm_group_bin_4145 (RW)
0x52: frame_vm_group_bin_20240 (RW)
0x53: frame_vm_group_bin_13044 (RW)
0x54: frame_vm_group_bin_19293 (RW)
0x55: frame_vm_group_bin_22059 (RW)
0x56: frame_vm_group_bin_14903 (RW)
0x57: frame_vm_group_bin_7688 (RW)
0x58: frame_vm_group_bin_13569 (RW)
0x59: frame_vm_group_bin_16718 (RW)
0x5: frame_vm_group_bin_12843 (RW)
0x5a: frame_vm_group_bin_9510 (RW)
0x5b: frame_vm_group_bin_2350 (RW)
0x5c: frame_vm_group_bin_18451 (RW)
0x5d: frame_vm_group_bin_11363 (RW)
0x5e: frame_vm_group_bin_4178 (RW)
0x5f: frame_vm_group_bin_20273 (RW)
0x60: frame_vm_group_bin_13078 (RW)
0x61: frame_vm_group_bin_0666 (RW)
0x62: frame_vm_group_bin_22088 (RW)
0x63: frame_vm_group_bin_14937 (RW)
0x64: frame_vm_group_bin_7721 (RW)
0x65: frame_vm_group_bin_18214 (RW)
0x66: frame_vm_group_bin_16752 (RW)
0x67: frame_vm_group_bin_9543 (RW)
0x68: frame_vm_group_bin_2383 (RW)
0x69: frame_vm_group_bin_18479 (RW)
0x6: frame_vm_group_bin_5769 (RW)
0x6a: frame_vm_group_bin_11395 (RW)
0x6b: frame_vm_group_bin_4210 (RW)
0x6c: frame_vm_group_bin_20306 (RW)
0x6d: frame_vm_group_bin_13111 (RW)
0x6e: frame_vm_group_bin_5961 (RW)
0x6f: frame_vm_group_bin_22119 (RW)
0x70: frame_vm_group_bin_14970 (RW)
0x71: frame_vm_group_bin_7754 (RW)
0x72: frame_vm_group_bin_0590 (RW)
0x73: frame_vm_group_bin_16785 (RW)
0x74: frame_vm_group_bin_9576 (RW)
0x75: frame_vm_group_bin_2416 (RW)
0x76: frame_vm_group_bin_18506 (RW)
0x77: frame_vm_group_bin_11427 (RW)
0x78: frame_vm_group_bin_4243 (RW)
0x79: frame_vm_group_bin_20341 (RW)
0x7: frame_vm_group_bin_21880 (RW)
0x7a: frame_vm_group_bin_13145 (RW)
0x7b: frame_vm_group_bin_5991 (RW)
0x7c: frame_vm_group_bin_22153 (RW)
0x7d: frame_vm_group_bin_15004 (RW)
0x7e: frame_vm_group_bin_7788 (RW)
0x7f: frame_vm_group_bin_4317 (RW)
0x80: frame_vm_group_bin_16819 (RW)
0x81: frame_vm_group_bin_9610 (RW)
0x82: frame_vm_group_bin_2449 (RW)
0x83: frame_vm_group_bin_18535 (RW)
0x84: frame_vm_group_bin_11461 (RW)
0x85: frame_vm_group_bin_4277 (RW)
0x86: frame_vm_group_bin_20375 (RW)
0x87: frame_vm_group_bin_13178 (RW)
0x88: frame_vm_group_bin_6021 (RW)
0x89: frame_vm_group_bin_22186 (RW)
0x8: frame_vm_group_bin_14705 (RW)
0x8a: frame_vm_group_bin_15035 (RW)
0x8b: frame_vm_group_bin_7821 (RW)
0x8c: frame_vm_group_bin_0656 (RW)
0x8d: frame_vm_group_bin_16852 (RW)
0x8e: frame_vm_group_bin_9643 (RW)
0x8f: frame_vm_group_bin_2481 (RW)
0x90: frame_vm_group_bin_18560 (RW)
0x91: frame_vm_group_bin_11494 (RW)
0x92: frame_vm_group_bin_4310 (RW)
0x93: frame_vm_group_bin_20408 (RW)
0x94: frame_vm_group_bin_13211 (RW)
0x95: frame_vm_group_bin_19317 (RW)
0x96: frame_vm_group_bin_22219 (RW)
0x97: frame_vm_group_bin_15060 (RW)
0x98: frame_vm_group_bin_7853 (RW)
0x99: frame_vm_group_bin_0689 (RW)
0x9: frame_vm_group_bin_7491 (RW)
0x9a: frame_vm_group_bin_16885 (RW)
0x9b: frame_vm_group_bin_9677 (RW)
0x9c: frame_vm_group_bin_2515 (RW)
0x9d: frame_vm_group_bin_18592 (RW)
0x9e: frame_vm_group_bin_11528 (RW)
0x9f: frame_vm_group_bin_4346 (RW)
0xa0: frame_vm_group_bin_20442 (RW)
0xa1: frame_vm_group_bin_13245 (RW)
0xa2: frame_vm_group_bin_0690 (RW)
0xa3: frame_vm_group_bin_22253 (RW)
0xa4: frame_vm_group_bin_15087 (RW)
0xa5: frame_vm_group_bin_7887 (RW)
0xa6: frame_vm_group_bin_0723 (RW)
0xa7: frame_vm_group_bin_16917 (RW)
0xa8: frame_vm_group_bin_9709 (RW)
0xa9: frame_vm_group_bin_2548 (RW)
0xa: frame_vm_group_bin_0337 (RW)
0xaa: frame_vm_group_bin_18625 (RW)
0xab: frame_vm_group_bin_11559 (RW)
0xac: frame_vm_group_bin_4379 (RW)
0xad: frame_vm_group_bin_20475 (RW)
0xae: frame_vm_group_bin_13278 (RW)
0xaf: frame_vm_group_bin_6104 (RW)
0xb0: frame_vm_group_bin_22285 (RW)
0xb1: frame_vm_group_bin_15111 (RW)
0xb2: frame_vm_group_bin_7920 (RW)
0xb3: frame_vm_group_bin_0756 (RW)
0xb4: frame_vm_group_bin_16950 (RW)
0xb5: frame_vm_group_bin_9742 (RW)
0xb6: frame_vm_group_bin_2581 (RW)
0xb7: frame_vm_group_bin_18657 (RW)
0xb8: frame_vm_group_bin_11586 (RW)
0xb9: frame_vm_group_bin_4412 (RW)
0xb: frame_vm_group_bin_16520 (RW)
0xba: frame_vm_group_bin_20509 (RW)
0xbb: frame_vm_group_bin_13312 (RW)
0xbc: frame_vm_group_bin_6137 (RW)
0xbd: frame_vm_group_bin_22319 (RW)
0xbe: frame_vm_group_bin_15138 (RW)
0xbf: frame_vm_group_bin_7955 (RW)
0xc0: frame_vm_group_bin_0790 (RW)
0xc1: frame_vm_group_bin_16984 (RW)
0xc2: frame_vm_group_bin_9776 (RW)
0xc3: frame_vm_group_bin_2615 (RW)
0xc4: frame_vm_group_bin_18691 (RW)
0xc5: frame_vm_group_bin_11614 (RW)
0xc6: frame_vm_group_bin_4446 (RW)
0xc7: frame_vm_group_bin_20542 (RW)
0xc8: frame_vm_group_bin_13344 (RW)
0xc9: frame_vm_group_bin_6169 (RW)
0xc: frame_vm_group_bin_9309 (RW)
0xca: frame_vm_group_bin_22351 (RW)
0xcb: frame_vm_group_bin_15167 (RW)
0xcc: frame_vm_group_bin_7987 (RW)
0xcd: frame_vm_group_bin_0822 (RW)
0xce: frame_vm_group_bin_17017 (RW)
0xcf: frame_vm_group_bin_9809 (RW)
0xd0: frame_vm_group_bin_2648 (RW)
0xd1: frame_vm_group_bin_18723 (RW)
0xd2: frame_vm_group_bin_1789 (RW)
0xd3: frame_vm_group_bin_4479 (RW)
0xd4: frame_vm_group_bin_20575 (RW)
0xd5: frame_vm_group_bin_13376 (RW)
0xd6: frame_vm_group_bin_6200 (RW)
0xd7: frame_vm_group_bin_22384 (RW)
0xd8: frame_vm_group_bin_15200 (RW)
0xd9: frame_vm_group_bin_8017 (RW)
0xd: frame_vm_group_bin_2158 (RW)
0xda: frame_vm_group_bin_0856 (RW)
0xdb: frame_vm_group_bin_17051 (RW)
0xdc: frame_vm_group_bin_9843 (RW)
0xdd: frame_vm_group_bin_2682 (RW)
0xde: frame_vm_group_bin_18755 (RW)
0xdf: frame_vm_group_bin_6426 (RW)
0xe0: frame_vm_group_bin_4513 (RW)
0xe1: frame_vm_group_bin_20609 (RW)
0xe2: frame_vm_group_bin_13409 (RW)
0xe3: frame_vm_group_bin_0713 (RW)
0xe4: frame_vm_group_bin_22417 (RW)
0xe5: frame_vm_group_bin_15235 (RW)
0xe6: frame_vm_group_bin_8047 (RW)
0xe7: frame_vm_group_bin_0889 (RW)
0xe8: frame_vm_group_bin_17084 (RW)
0xe9: frame_vm_group_bin_9876 (RW)
0xe: frame_vm_group_bin_18252 (RW)
0xea: frame_vm_group_bin_2715 (RW)
0xeb: frame_vm_group_bin_18788 (RW)
0xec: frame_vm_group_bin_11171 (RW)
0xed: frame_vm_group_bin_4546 (RW)
0xee: frame_vm_group_bin_20642 (RW)
0xef: frame_vm_group_bin_13442 (RW)
0xf0: frame_vm_group_bin_6258 (RW)
0xf1: frame_vm_group_bin_22450 (RW)
0xf2: frame_vm_group_bin_15268 (RW)
0xf3: frame_vm_group_bin_8078 (RW)
0xf4: frame_vm_group_bin_0922 (RW)
0xf5: frame_vm_group_bin_17117 (RW)
0xf6: frame_vm_group_bin_9908 (RW)
0xf7: frame_vm_group_bin_2748 (RW)
0xf8: frame_vm_group_bin_18821 (RW)
0xf9: frame_vm_group_bin_11710 (RW)
0xf: frame_vm_group_bin_11164 (RW)
0xfa: frame_vm_group_bin_4575 (RW)
0xfb: frame_vm_group_bin_20675 (RW)
0xfc: frame_vm_group_bin_13476 (RW)
0xfd: frame_vm_group_bin_6291 (RW)
0xfe: frame_vm_group_bin_22484 (RW)
0xff: frame_vm_group_bin_15301 (RW)
}
pt_vm_group_bin_0403 {
0x0: frame_vm_group_bin_3969 (RW)
0x100: frame_vm_group_bin_9963 (RW)
0x101: frame_vm_group_bin_2805 (RW)
0x102: frame_vm_group_bin_18879 (RW)
0x103: frame_vm_group_bin_11751 (RW)
0x104: frame_vm_group_bin_4615 (RW)
0x105: frame_vm_group_bin_20731 (RW)
0x106: frame_vm_group_bin_13532 (RW)
0x107: frame_vm_group_bin_6346 (RW)
0x108: frame_vm_group_bin_22539 (RW)
0x109: frame_vm_group_bin_15357 (RW)
0x10: frame_vm_group_bin_5807 (RW)
0x10a: frame_vm_group_bin_8166 (RW)
0x10b: frame_vm_group_bin_1011 (RW)
0x10c: frame_vm_group_bin_17203 (RW)
0x10d: frame_vm_group_bin_9996 (RW)
0x10e: frame_vm_group_bin_2838 (RW)
0x10f: frame_vm_group_bin_18912 (RW)
0x110: frame_vm_group_bin_11774 (RW)
0x111: frame_vm_group_bin_4643 (RW)
0x112: frame_vm_group_bin_20764 (RW)
0x113: frame_vm_group_bin_13565 (RW)
0x114: frame_vm_group_bin_6378 (RW)
0x115: frame_vm_group_bin_22572 (RW)
0x116: frame_vm_group_bin_15390 (RW)
0x117: frame_vm_group_bin_8199 (RW)
0x118: frame_vm_group_bin_1035 (RW)
0x119: frame_vm_group_bin_17235 (RW)
0x11: frame_vm_group_bin_21935 (RW)
0x11a: frame_vm_group_bin_10030 (RW)
0x11b: frame_vm_group_bin_2873 (RW)
0x11c: frame_vm_group_bin_18945 (RW)
0x11d: frame_vm_group_bin_11802 (RW)
0x11e: frame_vm_group_bin_4676 (RW)
0x11f: frame_vm_group_bin_20798 (RW)
0x120: frame_vm_group_bin_13599 (RW)
0x121: frame_vm_group_bin_6409 (RW)
0x122: frame_vm_group_bin_22606 (RW)
0x123: frame_vm_group_bin_15424 (RW)
0x124: frame_vm_group_bin_8233 (RW)
0x125: frame_vm_group_bin_1057 (RW)
0x126: frame_vm_group_bin_17269 (RW)
0x127: frame_vm_group_bin_10063 (RW)
0x128: frame_vm_group_bin_2906 (RW)
0x129: frame_vm_group_bin_18976 (RW)
0x12: frame_vm_group_bin_14760 (RW)
0x12a: frame_vm_group_bin_11835 (RW)
0x12b: frame_vm_group_bin_4708 (RW)
0x12c: frame_vm_group_bin_20830 (RW)
0x12d: frame_vm_group_bin_13632 (RW)
0x12e: frame_vm_group_bin_6442 (RW)
0x12f: frame_vm_group_bin_22639 (RW)
0x130: frame_vm_group_bin_15457 (RW)
0x131: frame_vm_group_bin_8266 (RW)
0x132: frame_vm_group_bin_1081 (RW)
0x133: frame_vm_group_bin_17302 (RW)
0x134: frame_vm_group_bin_10096 (RW)
0x135: frame_vm_group_bin_2939 (RW)
0x136: frame_vm_group_bin_19009 (RW)
0x137: frame_vm_group_bin_11863 (RW)
0x138: frame_vm_group_bin_4740 (RW)
0x139: frame_vm_group_bin_20858 (RW)
0x13: frame_vm_group_bin_7545 (RW)
0x13a: frame_vm_group_bin_13665 (RW)
0x13b: frame_vm_group_bin_6476 (RW)
0x13c: frame_vm_group_bin_22673 (RW)
0x13d: frame_vm_group_bin_15491 (RW)
0x13e: frame_vm_group_bin_8299 (RW)
0x13f: frame_vm_group_bin_1111 (RW)
0x140: frame_vm_group_bin_17336 (RW)
0x141: frame_vm_group_bin_10130 (RW)
0x142: frame_vm_group_bin_2973 (RW)
0x143: frame_vm_group_bin_19043 (RW)
0x144: frame_vm_group_bin_11891 (RW)
0x145: frame_vm_group_bin_4774 (RW)
0x146: frame_vm_group_bin_20883 (RW)
0x147: frame_vm_group_bin_13698 (RW)
0x148: frame_vm_group_bin_6509 (RW)
0x149: frame_vm_group_bin_22706 (RW)
0x14: frame_vm_group_bin_0390 (RW)
0x14a: frame_vm_group_bin_15523 (RW)
0x14b: frame_vm_group_bin_8332 (RW)
0x14c: frame_vm_group_bin_1143 (RW)
0x14d: frame_vm_group_bin_17368 (RW)
0x14e: frame_vm_group_bin_10165 (RW)
0x14f: frame_vm_group_bin_3006 (RW)
0x150: frame_vm_group_bin_19076 (RW)
0x151: frame_vm_group_bin_11915 (RW)
0x152: frame_vm_group_bin_4807 (RW)
0x153: frame_vm_group_bin_20911 (RW)
0x154: frame_vm_group_bin_13730 (RW)
0x155: frame_vm_group_bin_6542 (RW)
0x156: frame_vm_group_bin_22739 (RW)
0x157: frame_vm_group_bin_15555 (RW)
0x158: frame_vm_group_bin_8365 (RW)
0x159: frame_vm_group_bin_1176 (RW)
0x15: frame_vm_group_bin_16575 (RW)
0x15a: frame_vm_group_bin_17399 (RW)
0x15b: frame_vm_group_bin_10199 (RW)
0x15c: frame_vm_group_bin_3040 (RW)
0x15d: frame_vm_group_bin_19109 (RW)
0x15e: frame_vm_group_bin_11945 (RW)
0x15f: frame_vm_group_bin_4840 (RW)
0x160: frame_vm_group_bin_20941 (RW)
0x161: frame_vm_group_bin_13765 (RW)
0x162: frame_vm_group_bin_6576 (RW)
0x163: frame_vm_group_bin_22772 (RW)
0x164: frame_vm_group_bin_15589 (RW)
0x165: frame_vm_group_bin_8399 (RW)
0x166: frame_vm_group_bin_1210 (RW)
0x167: frame_vm_group_bin_17424 (RW)
0x168: frame_vm_group_bin_10232 (RW)
0x169: frame_vm_group_bin_3073 (RW)
0x16: frame_vm_group_bin_9364 (RW)
0x16a: frame_vm_group_bin_19141 (RW)
0x16b: frame_vm_group_bin_11978 (RW)
0x16c: frame_vm_group_bin_4873 (RW)
0x16d: frame_vm_group_bin_20966 (RW)
0x16e: frame_vm_group_bin_13798 (RW)
0x16f: frame_vm_group_bin_6609 (RW)
0x170: frame_vm_group_bin_22805 (RW)
0x171: frame_vm_group_bin_15622 (RW)
0x172: frame_vm_group_bin_8432 (RW)
0x173: frame_vm_group_bin_1243 (RW)
0x174: frame_vm_group_bin_17449 (RW)
0x175: frame_vm_group_bin_10265 (RW)
0x176: frame_vm_group_bin_3106 (RW)
0x177: frame_vm_group_bin_19174 (RW)
0x178: frame_vm_group_bin_12010 (RW)
0x179: frame_vm_group_bin_4906 (RW)
0x17: frame_vm_group_bin_2210 (RW)
0x17a: frame_vm_group_bin_21000 (RW)
0x17b: frame_vm_group_bin_13830 (RW)
0x17c: frame_vm_group_bin_6643 (RW)
0x17d: frame_vm_group_bin_22839 (RW)
0x17e: frame_vm_group_bin_15656 (RW)
0x17f: frame_vm_group_bin_8466 (RW)
0x180: frame_vm_group_bin_1274 (RW)
0x181: frame_vm_group_bin_17470 (RW)
0x182: frame_vm_group_bin_10299 (RW)
0x183: frame_vm_group_bin_3139 (RW)
0x184: frame_vm_group_bin_19208 (RW)
0x185: frame_vm_group_bin_12041 (RW)
0x186: frame_vm_group_bin_4938 (RW)
0x187: frame_vm_group_bin_21033 (RW)
0x188: frame_vm_group_bin_13859 (RW)
0x189: frame_vm_group_bin_6676 (RW)
0x18: frame_vm_group_bin_18308 (RW)
0x18a: frame_vm_group_bin_22872 (RW)
0x18b: frame_vm_group_bin_15689 (RW)
0x18c: frame_vm_group_bin_8499 (RW)
0x18d: frame_vm_group_bin_1307 (RW)
0x18e: frame_vm_group_bin_17492 (RW)
0x18f: frame_vm_group_bin_10332 (RW)
0x190: frame_vm_group_bin_3172 (RW)
0x191: frame_vm_group_bin_19241 (RW)
0x192: frame_vm_group_bin_12068 (RW)
0x193: frame_vm_group_bin_4969 (RW)
0x194: frame_vm_group_bin_21067 (RW)
0x195: frame_vm_group_bin_13889 (RW)
0x196: frame_vm_group_bin_6709 (RW)
0x197: frame_vm_group_bin_22905 (RW)
0x198: frame_vm_group_bin_15722 (RW)
0x199: frame_vm_group_bin_8531 (RW)
0x19: frame_vm_group_bin_11220 (RW)
0x19a: frame_vm_group_bin_1340 (RW)
0x19b: frame_vm_group_bin_17518 (RW)
0x19c: frame_vm_group_bin_10366 (RW)
0x19d: frame_vm_group_bin_3206 (RW)
0x19e: frame_vm_group_bin_19275 (RW)
0x19f: frame_vm_group_bin_12102 (RW)
0x1: frame_vm_group_bin_20066 (RW)
0x1a0: frame_vm_group_bin_5003 (RW)
0x1a1: frame_vm_group_bin_21101 (RW)
0x1a2: frame_vm_group_bin_13923 (RW)
0x1a3: frame_vm_group_bin_6742 (RW)
0x1a4: frame_vm_group_bin_22939 (RW)
0x1a5: frame_vm_group_bin_15756 (RW)
0x1a6: frame_vm_group_bin_8563 (RW)
0x1a7: frame_vm_group_bin_1374 (RW)
0x1a8: frame_vm_group_bin_17544 (RW)
0x1a9: frame_vm_group_bin_10395 (RW)
0x1a: frame_vm_group_bin_4036 (RW)
0x1aa: frame_vm_group_bin_3238 (RW)
0x1ab: frame_vm_group_bin_19308 (RW)
0x1ac: frame_vm_group_bin_12134 (RW)
0x1ad: frame_vm_group_bin_5036 (RW)
0x1ae: frame_vm_group_bin_21134 (RW)
0x1af: frame_vm_group_bin_13956 (RW)
0x1b0: frame_vm_group_bin_6774 (RW)
0x1b1: frame_vm_group_bin_22971 (RW)
0x1b2: frame_vm_group_bin_15789 (RW)
0x1b3: frame_vm_group_bin_8596 (RW)
0x1b4: frame_vm_group_bin_1407 (RW)
0x1b5: frame_vm_group_bin_17565 (RW)
0x1b6: frame_vm_group_bin_10421 (RW)
0x1b7: frame_vm_group_bin_3271 (RW)
0x1b8: frame_vm_group_bin_19341 (RW)
0x1b9: frame_vm_group_bin_12165 (RW)
0x1b: frame_vm_group_bin_20132 (RW)
0x1ba: frame_vm_group_bin_5071 (RW)
0x1bb: frame_vm_group_bin_21167 (RW)
0x1bc: frame_vm_group_bin_13990 (RW)
0x1bd: frame_vm_group_bin_6808 (RW)
0x1be: frame_vm_group_bin_23004 (RW)
0x1bf: frame_vm_group_bin_15821 (RW)
0x1c0: frame_vm_group_bin_8629 (RW)
0x1c1: frame_vm_group_bin_1441 (RW)
0x1c2: frame_vm_group_bin_17590 (RW)
0x1c3: frame_vm_group_bin_10452 (RW)
0x1c4: frame_vm_group_bin_3305 (RW)
0x1c5: frame_vm_group_bin_19375 (RW)
0x1c6: frame_vm_group_bin_12197 (RW)
0x1c7: frame_vm_group_bin_5104 (RW)
0x1c8: frame_vm_group_bin_21200 (RW)
0x1c9: frame_vm_group_bin_14023 (RW)
0x1c: frame_vm_group_bin_12932 (RW)
0x1ca: frame_vm_group_bin_6836 (RW)
0x1cb: frame_vm_group_bin_23037 (RW)
0x1cc: frame_vm_group_bin_15854 (RW)
0x1cd: frame_vm_group_bin_8662 (RW)
0x1ce: frame_vm_group_bin_1474 (RW)
0x1cf: frame_vm_group_bin_17614 (RW)
0x1d0: frame_vm_group_bin_10485 (RW)
0x1d1: frame_vm_group_bin_3338 (RW)
0x1d2: frame_vm_group_bin_19408 (RW)
0x1d3: frame_vm_group_bin_12227 (RW)
0x1d4: frame_vm_group_bin_5137 (RW)
0x1d5: frame_vm_group_bin_21233 (RW)
0x1d6: frame_vm_group_bin_14056 (RW)
0x1d7: frame_vm_group_bin_6863 (RW)
0x1d8: frame_vm_group_bin_23070 (RW)
0x1d9: frame_vm_group_bin_15887 (RW)
0x1d: frame_vm_group_bin_5830 (RW)
0x1da: frame_vm_group_bin_8697 (RW)
0x1db: frame_vm_group_bin_1508 (RW)
0x1dc: frame_vm_group_bin_17648 (RW)
0x1dd: frame_vm_group_bin_10518 (RW)
0x1de: frame_vm_group_bin_3372 (RW)
0x1df: frame_vm_group_bin_19439 (RW)
0x1e0: frame_vm_group_bin_12260 (RW)
0x1e1: frame_vm_group_bin_5171 (RW)
0x1e2: frame_vm_group_bin_21267 (RW)
0x1e3: frame_vm_group_bin_14090 (RW)
0x1e4: frame_vm_group_bin_6889 (RW)
0x1e5: frame_vm_group_bin_23104 (RW)
0x1e6: frame_vm_group_bin_15921 (RW)
0x1e7: frame_vm_group_bin_8730 (RW)
0x1e8: frame_vm_group_bin_1541 (RW)
0x1e9: frame_vm_group_bin_17681 (RW)
0x1e: frame_vm_group_bin_21969 (RW)
0x1ea: frame_vm_group_bin_10551 (RW)
0x1eb: frame_vm_group_bin_3400 (RW)
0x1ec: frame_vm_group_bin_19471 (RW)
0x1ed: frame_vm_group_bin_12293 (RW)
0x1ee: frame_vm_group_bin_5204 (RW)
0x1ef: frame_vm_group_bin_21300 (RW)
0x1f0: frame_vm_group_bin_14123 (RW)
0x1f1: frame_vm_group_bin_6913 (RW)
0x1f2: frame_vm_group_bin_23137 (RW)
0x1f3: frame_vm_group_bin_15954 (RW)
0x1f4: frame_vm_group_bin_8763 (RW)
0x1f5: frame_vm_group_bin_1574 (RW)
0x1f6: frame_vm_group_bin_17707 (RW)
0x1f7: frame_vm_group_bin_10584 (RW)
0x1f8: frame_vm_group_bin_3424 (RW)
0x1f9: frame_vm_group_bin_19504 (RW)
0x1f: frame_vm_group_bin_14793 (RW)
0x1fa: frame_vm_group_bin_12326 (RW)
0x1fb: frame_vm_group_bin_5238 (RW)
0x1fc: frame_vm_group_bin_21332 (RW)
0x1fd: frame_vm_group_bin_14157 (RW)
0x1fe: frame_vm_group_bin_6944 (RW)
0x1ff: frame_vm_group_bin_23170 (RW)
0x20: frame_vm_group_bin_7578 (RW)
0x21: frame_vm_group_bin_0419 (RW)
0x22: frame_vm_group_bin_16608 (RW)
0x23: frame_vm_group_bin_9399 (RW)
0x24: frame_vm_group_bin_2240 (RW)
0x25: frame_vm_group_bin_18342 (RW)
0x26: frame_vm_group_bin_11254 (RW)
0x27: frame_vm_group_bin_4069 (RW)
0x28: frame_vm_group_bin_20164 (RW)
0x29: frame_vm_group_bin_12965 (RW)
0x2: frame_vm_group_bin_12866 (RW)
0x2a: frame_vm_group_bin_5854 (RW)
0x2b: frame_vm_group_bin_22002 (RW)
0x2c: frame_vm_group_bin_14826 (RW)
0x2d: frame_vm_group_bin_7611 (RW)
0x2e: frame_vm_group_bin_0451 (RW)
0x2f: frame_vm_group_bin_16641 (RW)
0x30: frame_vm_group_bin_9432 (RW)
0x31: frame_vm_group_bin_2272 (RW)
0x32: frame_vm_group_bin_18375 (RW)
0x33: frame_vm_group_bin_11287 (RW)
0x34: frame_vm_group_bin_4102 (RW)
0x35: frame_vm_group_bin_20196 (RW)
0x36: frame_vm_group_bin_12998 (RW)
0x37: frame_vm_group_bin_5880 (RW)
0x38: frame_vm_group_bin_22029 (RW)
0x39: frame_vm_group_bin_14859 (RW)
0x3: frame_vm_group_bin_5785 (RW)
0x3a: frame_vm_group_bin_7645 (RW)
0x3b: frame_vm_group_bin_0484 (RW)
0x3c: frame_vm_group_bin_16675 (RW)
0x3d: frame_vm_group_bin_9466 (RW)
0x3e: frame_vm_group_bin_2306 (RW)
0x3f: frame_vm_group_bin_18407 (RW)
0x40: frame_vm_group_bin_11321 (RW)
0x41: frame_vm_group_bin_4135 (RW)
0x42: frame_vm_group_bin_20230 (RW)
0x43: frame_vm_group_bin_13034 (RW)
0x44: frame_vm_group_bin_5907 (RW)
0x45: frame_vm_group_bin_22051 (RW)
0x46: frame_vm_group_bin_14893 (RW)
0x47: frame_vm_group_bin_7678 (RW)
0x48: frame_vm_group_bin_0517 (RW)
0x49: frame_vm_group_bin_16707 (RW)
0x4: frame_vm_group_bin_21903 (RW)
0x4a: frame_vm_group_bin_9499 (RW)
0x4b: frame_vm_group_bin_2339 (RW)
0x4c: frame_vm_group_bin_18440 (RW)
0x4d: frame_vm_group_bin_11352 (RW)
0x4e: frame_vm_group_bin_4167 (RW)
0x4f: frame_vm_group_bin_20263 (RW)
0x50: frame_vm_group_bin_13067 (RW)
0x51: frame_vm_group_bin_5932 (RW)
0x52: frame_vm_group_bin_22077 (RW)
0x53: frame_vm_group_bin_14926 (RW)
0x54: frame_vm_group_bin_7711 (RW)
0x55: frame_vm_group_bin_0549 (RW)
0x56: frame_vm_group_bin_16741 (RW)
0x57: frame_vm_group_bin_9532 (RW)
0x58: frame_vm_group_bin_2372 (RW)
0x59: frame_vm_group_bin_18471 (RW)
0x5: frame_vm_group_bin_14728 (RW)
0x5a: frame_vm_group_bin_11385 (RW)
0x5b: frame_vm_group_bin_4200 (RW)
0x5c: frame_vm_group_bin_20296 (RW)
0x5d: frame_vm_group_bin_13101 (RW)
0x5e: frame_vm_group_bin_5954 (RW)
0x5f: frame_vm_group_bin_22109 (RW)
0x60: frame_vm_group_bin_14960 (RW)
0x61: frame_vm_group_bin_7744 (RW)
0x62: frame_vm_group_bin_0581 (RW)
0x63: frame_vm_group_bin_16775 (RW)
0x64: frame_vm_group_bin_9566 (RW)
0x65: frame_vm_group_bin_2406 (RW)
0x66: frame_vm_group_bin_18498 (RW)
0x67: frame_vm_group_bin_11417 (RW)
0x68: frame_vm_group_bin_4233 (RW)
0x69: frame_vm_group_bin_20331 (RW)
0x6: frame_vm_group_bin_7513 (RW)
0x6a: frame_vm_group_bin_13134 (RW)
0x6b: frame_vm_group_bin_5981 (RW)
0x6c: frame_vm_group_bin_22142 (RW)
0x6d: frame_vm_group_bin_14993 (RW)
0x6e: frame_vm_group_bin_7777 (RW)
0x6f: frame_vm_group_bin_0613 (RW)
0x70: frame_vm_group_bin_16808 (RW)
0x71: frame_vm_group_bin_9599 (RW)
0x72: frame_vm_group_bin_2438 (RW)
0x73: frame_vm_group_bin_18524 (RW)
0x74: frame_vm_group_bin_11450 (RW)
0x75: frame_vm_group_bin_4266 (RW)
0x76: frame_vm_group_bin_20364 (RW)
0x77: frame_vm_group_bin_13167 (RW)
0x78: frame_vm_group_bin_6012 (RW)
0x79: frame_vm_group_bin_22175 (RW)
0x7: frame_vm_group_bin_0359 (RW)
0x7a: frame_vm_group_bin_15027 (RW)
0x7b: frame_vm_group_bin_7811 (RW)
0x7c: frame_vm_group_bin_0646 (RW)
0x7d: frame_vm_group_bin_16842 (RW)
0x7e: frame_vm_group_bin_9633 (RW)
0x7f: frame_vm_group_bin_2471 (RW)
0x80: frame_vm_group_bin_18552 (RW)
0x81: frame_vm_group_bin_11484 (RW)
0x82: frame_vm_group_bin_4300 (RW)
0x83: frame_vm_group_bin_20398 (RW)
0x84: frame_vm_group_bin_13201 (RW)
0x85: frame_vm_group_bin_6043 (RW)
0x86: frame_vm_group_bin_22209 (RW)
0x87: frame_vm_group_bin_15052 (RW)
0x88: frame_vm_group_bin_7843 (RW)
0x89: frame_vm_group_bin_0679 (RW)
0x8: frame_vm_group_bin_16543 (RW)
0x8a: frame_vm_group_bin_16874 (RW)
0x8b: frame_vm_group_bin_9666 (RW)
0x8c: frame_vm_group_bin_2504 (RW)
0x8d: frame_vm_group_bin_18581 (RW)
0x8e: frame_vm_group_bin_11517 (RW)
0x8f: frame_vm_group_bin_4333 (RW)
0x90: frame_vm_group_bin_20431 (RW)
0x91: frame_vm_group_bin_13234 (RW)
0x92: frame_vm_group_bin_6066 (RW)
0x93: frame_vm_group_bin_22242 (RW)
0x94: frame_vm_group_bin_15076 (RW)
0x95: frame_vm_group_bin_7876 (RW)
0x96: frame_vm_group_bin_0712 (RW)
0x97: frame_vm_group_bin_16906 (RW)
0x98: frame_vm_group_bin_9698 (RW)
0x99: frame_vm_group_bin_2537 (RW)
0x9: frame_vm_group_bin_9331 (RW)
0x9a: frame_vm_group_bin_18615 (RW)
0x9b: frame_vm_group_bin_11551 (RW)
0x9c: frame_vm_group_bin_4369 (RW)
0x9d: frame_vm_group_bin_20465 (RW)
0x9e: frame_vm_group_bin_13268 (RW)
0x9f: frame_vm_group_bin_6095 (RW)
0xa0: frame_vm_group_bin_22275 (RW)
0xa1: frame_vm_group_bin_15104 (RW)
0xa2: frame_vm_group_bin_7910 (RW)
0xa3: frame_vm_group_bin_0746 (RW)
0xa4: frame_vm_group_bin_16940 (RW)
0xa5: frame_vm_group_bin_9732 (RW)
0xa6: frame_vm_group_bin_2571 (RW)
0xa7: frame_vm_group_bin_18647 (RW)
0xa8: frame_vm_group_bin_11579 (RW)
0xa9: frame_vm_group_bin_4402 (RW)
0xa: frame_vm_group_bin_2181 (RW)
0xaa: frame_vm_group_bin_20498 (RW)
0xab: frame_vm_group_bin_13301 (RW)
0xac: frame_vm_group_bin_6126 (RW)
0xad: frame_vm_group_bin_22308 (RW)
0xae: frame_vm_group_bin_15130 (RW)
0xaf: frame_vm_group_bin_7944 (RW)
0xb0: frame_vm_group_bin_0779 (RW)
0xb1: frame_vm_group_bin_16973 (RW)
0xb2: frame_vm_group_bin_9765 (RW)
0xb3: frame_vm_group_bin_2604 (RW)
0xb4: frame_vm_group_bin_18680 (RW)
0xb5: frame_vm_group_bin_11603 (RW)
0xb6: frame_vm_group_bin_4435 (RW)
0xb7: frame_vm_group_bin_20531 (RW)
0xb8: frame_vm_group_bin_13333 (RW)
0xb9: frame_vm_group_bin_6158 (RW)
0xb: frame_vm_group_bin_18275 (RW)
0xba: frame_vm_group_bin_22341 (RW)
0xbb: frame_vm_group_bin_15157 (RW)
0xbc: frame_vm_group_bin_7978 (RW)
0xbd: frame_vm_group_bin_0812 (RW)
0xbe: frame_vm_group_bin_17007 (RW)
0xbf: frame_vm_group_bin_9799 (RW)
0xc0: frame_vm_group_bin_2638 (RW)
0xc1: frame_vm_group_bin_18713 (RW)
0xc2: frame_vm_group_bin_11631 (RW)
0xc3: frame_vm_group_bin_4469 (RW)
0xc4: frame_vm_group_bin_20565 (RW)
0xc5: frame_vm_group_bin_13367 (RW)
0xc6: frame_vm_group_bin_6191 (RW)
0xc7: frame_vm_group_bin_22374 (RW)
0xc8: frame_vm_group_bin_15190 (RW)
0xc9: frame_vm_group_bin_8008 (RW)
0xc: frame_vm_group_bin_11187 (RW)
0xca: frame_vm_group_bin_0845 (RW)
0xcb: frame_vm_group_bin_17040 (RW)
0xcc: frame_vm_group_bin_9832 (RW)
0xcd: frame_vm_group_bin_2671 (RW)
0xce: frame_vm_group_bin_18744 (RW)
0xcf: frame_vm_group_bin_11653 (RW)
0xd0: frame_vm_group_bin_4502 (RW)
0xd1: frame_vm_group_bin_20598 (RW)
0xd2: frame_vm_group_bin_13398 (RW)
0xd3: frame_vm_group_bin_6218 (RW)
0xd4: frame_vm_group_bin_22407 (RW)
0xd5: frame_vm_group_bin_15223 (RW)
0xd6: frame_vm_group_bin_8036 (RW)
0xd7: frame_vm_group_bin_0878 (RW)
0xd8: frame_vm_group_bin_17073 (RW)
0xd9: frame_vm_group_bin_9865 (RW)
0xd: frame_vm_group_bin_4002 (RW)
0xda: frame_vm_group_bin_2705 (RW)
0xdb: frame_vm_group_bin_18778 (RW)
0xdc: frame_vm_group_bin_11674 (RW)
0xdd: frame_vm_group_bin_4536 (RW)
0xde: frame_vm_group_bin_20632 (RW)
0xdf: frame_vm_group_bin_13432 (RW)
0xe0: frame_vm_group_bin_6248 (RW)
0xe1: frame_vm_group_bin_22440 (RW)
0xe2: frame_vm_group_bin_15258 (RW)
0xe3: frame_vm_group_bin_8068 (RW)
0xe4: frame_vm_group_bin_0912 (RW)
0xe5: frame_vm_group_bin_17107 (RW)
0xe6: frame_vm_group_bin_9898 (RW)
0xe7: frame_vm_group_bin_2738 (RW)
0xe8: frame_vm_group_bin_18811 (RW)
0xe9: frame_vm_group_bin_11701 (RW)
0xe: frame_vm_group_bin_20099 (RW)
0xea: frame_vm_group_bin_4567 (RW)
0xeb: frame_vm_group_bin_20664 (RW)
0xec: frame_vm_group_bin_13465 (RW)
0xed: frame_vm_group_bin_6280 (RW)
0xee: frame_vm_group_bin_22473 (RW)
0xef: frame_vm_group_bin_15290 (RW)
0xf0: frame_vm_group_bin_8100 (RW)
0xf1: frame_vm_group_bin_0945 (RW)
0xf2: frame_vm_group_bin_17140 (RW)
0xf3: frame_vm_group_bin_9931 (RW)
0xf4: frame_vm_group_bin_2771 (RW)
0xf5: frame_vm_group_bin_18845 (RW)
0xf6: frame_vm_group_bin_11728 (RW)
0xf7: frame_vm_group_bin_4590 (RW)
0xf8: frame_vm_group_bin_20697 (RW)
0xf9: frame_vm_group_bin_13498 (RW)
0xf: frame_vm_group_bin_12899 (RW)
0xfa: frame_vm_group_bin_6314 (RW)
0xfb: frame_vm_group_bin_22507 (RW)
0xfc: frame_vm_group_bin_15324 (RW)
0xfd: frame_vm_group_bin_8133 (RW)
0xfe: frame_vm_group_bin_0979 (RW)
0xff: frame_vm_group_bin_17172 (RW)
}
pt_vm_group_bin_1120 {
0x0: frame_vm_group_bin_4700 (RW)
0x10: frame_vm_group_bin_6467 (RW)
0x11: frame_vm_group_bin_22664 (RW)
0x12: frame_vm_group_bin_15482 (RW)
0x13: frame_vm_group_bin_8290 (RW)
0x14: frame_vm_group_bin_1102 (RW)
0x15: frame_vm_group_bin_17327 (RW)
0x16: frame_vm_group_bin_10121 (RW)
0x17: frame_vm_group_bin_2964 (RW)
0x18: frame_vm_group_bin_19034 (RW)
0x19: frame_vm_group_bin_11885 (RW)
0x1: frame_vm_group_bin_20822 (RW)
0x1a: frame_vm_group_bin_4766 (RW)
0x1b: frame_vm_group_bin_20877 (RW)
0x1c: frame_vm_group_bin_13690 (RW)
0x1d: frame_vm_group_bin_6501 (RW)
0x1e: frame_vm_group_bin_22698 (RW)
0x1f: frame_vm_group_bin_15515 (RW)
0x20: frame_vm_group_bin_8324 (RW)
0x21: frame_vm_group_bin_1135 (RW)
0x22: frame_vm_group_bin_17360 (RW)
0x23: frame_vm_group_bin_10157 (RW)
0x24: frame_vm_group_bin_2998 (RW)
0x25: frame_vm_group_bin_19068 (RW)
0x26: frame_vm_group_bin_11909 (RW)
0x27: frame_vm_group_bin_4799 (RW)
0x28: frame_vm_group_bin_20904 (RW)
0x29: frame_vm_group_bin_13722 (RW)
0x2: frame_vm_group_bin_13624 (RW)
0x2a: frame_vm_group_bin_6534 (RW)
0x2b: frame_vm_group_bin_22731 (RW)
0x2c: frame_vm_group_bin_15547 (RW)
0x2d: frame_vm_group_bin_8357 (RW)
0x2e: frame_vm_group_bin_1168 (RW)
0x2f: frame_vm_group_bin_17390 (RW)
0x30: frame_vm_group_bin_10190 (RW)
0x31: frame_vm_group_bin_3031 (RW)
0x32: frame_vm_group_bin_19101 (RW)
0x33: frame_vm_group_bin_11939 (RW)
0x34: frame_vm_group_bin_4831 (RW)
0x35: frame_vm_group_bin_20932 (RW)
0x36: frame_vm_group_bin_13755 (RW)
0x37: frame_vm_group_bin_6567 (RW)
0x38: frame_vm_group_bin_22763 (RW)
0x39: frame_vm_group_bin_15580 (RW)
0x3: frame_vm_group_bin_6434 (RW)
0x3a: frame_vm_group_bin_8391 (RW)
0x3b: frame_vm_group_bin_1202 (RW)
0x3c: frame_vm_group_bin_17418 (RW)
0x3d: frame_vm_group_bin_10224 (RW)
0x3e: frame_vm_group_bin_3065 (RW)
0x3f: frame_vm_group_bin_19133 (RW)
0x40: frame_vm_group_bin_11970 (RW)
0x41: frame_vm_group_bin_4865 (RW)
0x42: frame_vm_group_bin_20960 (RW)
0x43: frame_vm_group_bin_13790 (RW)
0x44: frame_vm_group_bin_6601 (RW)
0x45: frame_vm_group_bin_22797 (RW)
0x46: frame_vm_group_bin_15614 (RW)
0x47: frame_vm_group_bin_8424 (RW)
0x48: frame_vm_group_bin_1235 (RW)
0x49: frame_vm_group_bin_17443 (RW)
0x4: frame_vm_group_bin_22631 (RW)
0x4a: frame_vm_group_bin_10257 (RW)
0x4b: frame_vm_group_bin_3098 (RW)
0x4c: frame_vm_group_bin_19166 (RW)
0x4d: frame_vm_group_bin_12002 (RW)
0x4e: frame_vm_group_bin_4898 (RW)
0x4f: frame_vm_group_bin_20991 (RW)
0x50: frame_vm_group_bin_13821 (RW)
0x51: frame_vm_group_bin_6634 (RW)
0x52: frame_vm_group_bin_22830 (RW)
0x53: frame_vm_group_bin_15647 (RW)
0x54: frame_vm_group_bin_8457 (RW)
0x55: frame_vm_group_bin_1267 (RW)
0x56: frame_vm_group_bin_17465 (RW)
0x57: frame_vm_group_bin_10290 (RW)
0x58: frame_vm_group_bin_3130 (RW)
0x59: frame_vm_group_bin_19199 (RW)
0x5: frame_vm_group_bin_15449 (RW)
0x5a: frame_vm_group_bin_12033 (RW)
0x5b: frame_vm_group_bin_4930 (RW)
0x5c: frame_vm_group_bin_21025 (RW)
0x5d: frame_vm_group_bin_13852 (RW)
0x5e: frame_vm_group_bin_6668 (RW)
0x5f: frame_vm_group_bin_22864 (RW)
0x60: frame_vm_group_bin_15681 (RW)
0x61: frame_vm_group_bin_8491 (RW)
0x62: frame_vm_group_bin_1299 (RW)
0x63: frame_vm_group_bin_17486 (RW)
0x64: frame_vm_group_bin_10324 (RW)
0x65: frame_vm_group_bin_3164 (RW)
0x66: frame_vm_group_bin_19233 (RW)
0x67: frame_vm_group_bin_12061 (RW)
0x68: frame_vm_group_bin_4962 (RW)
0x69: frame_vm_group_bin_21059 (RW)
0x6: frame_vm_group_bin_8258 (RW)
0x6a: frame_vm_group_bin_13881 (RW)
0x6b: frame_vm_group_bin_6701 (RW)
0x6c: frame_vm_group_bin_22897 (RW)
0x6d: frame_vm_group_bin_15714 (RW)
0x6e: frame_vm_group_bin_8523 (RW)
0x6f: frame_vm_group_bin_1331 (RW)
0x70: frame_vm_group_bin_17510 (RW)
0x71: frame_vm_group_bin_10357 (RW)
0x72: frame_vm_group_bin_3197 (RW)
0x73: frame_vm_group_bin_19266 (RW)
0x74: frame_vm_group_bin_12093 (RW)
0x75: frame_vm_group_bin_4994 (RW)
0x76: frame_vm_group_bin_21092 (RW)
0x77: frame_vm_group_bin_13914 (RW)
0x78: frame_vm_group_bin_6733 (RW)
0x79: frame_vm_group_bin_22930 (RW)
0x7: frame_vm_group_bin_1075 (RW)
0x7a: frame_vm_group_bin_15748 (RW)
0x7b: frame_vm_group_bin_8555 (RW)
0x7c: frame_vm_group_bin_1367 (RW)
0x7d: frame_vm_group_bin_17539 (RW)
0x7e: frame_vm_group_bin_10390 (RW)
0x7f: frame_vm_group_bin_3230 (RW)
0x80: frame_vm_group_bin_19300 (RW)
0x81: frame_vm_group_bin_12126 (RW)
0x82: frame_vm_group_bin_5028 (RW)
0x83: frame_vm_group_bin_21126 (RW)
0x84: frame_vm_group_bin_13948 (RW)
0x85: frame_vm_group_bin_6766 (RW)
0x86: frame_vm_group_bin_22963 (RW)
0x87: frame_vm_group_bin_15781 (RW)
0x88: frame_vm_group_bin_8588 (RW)
0x89: frame_vm_group_bin_1399 (RW)
0x8: frame_vm_group_bin_17294 (RW)
0x8a: frame_vm_group_bin_17560 (RW)
0x8b: frame_vm_group_bin_10415 (RW)
0x8c: frame_vm_group_bin_3263 (RW)
0x8d: frame_vm_group_bin_19333 (RW)
0x8e: frame_vm_group_bin_12159 (RW)
0x8f: frame_vm_group_bin_5061 (RW)
0x90: frame_vm_group_bin_21158 (RW)
0x91: frame_vm_group_bin_13981 (RW)
0x92: frame_vm_group_bin_6799 (RW)
0x93: frame_vm_group_bin_22996 (RW)
0x94: frame_vm_group_bin_15813 (RW)
0x95: frame_vm_group_bin_8620 (RW)
0x96: frame_vm_group_bin_1432 (RW)
0x97: frame_vm_group_bin_17583 (RW)
0x98: frame_vm_group_bin_10443 (RW)
0x99: frame_vm_group_bin_3296 (RW)
0x9: frame_vm_group_bin_10088 (RW)
0x9a: frame_vm_group_bin_19367 (RW)
0x9b: frame_vm_group_bin_12189 (RW)
0x9c: frame_vm_group_bin_5096 (RW)
0x9d: frame_vm_group_bin_21192 (RW)
0x9e: frame_vm_group_bin_14015 (RW)
0x9f: frame_vm_group_bin_6830 (RW)
0xa0: frame_vm_group_bin_23029 (RW)
0xa1: frame_vm_group_bin_15846 (RW)
0xa2: frame_vm_group_bin_8654 (RW)
0xa3: frame_vm_group_bin_1466 (RW)
0xa4: frame_vm_group_bin_17608 (RW)
0xa5: frame_vm_group_bin_10477 (RW)
0xa6: frame_vm_group_bin_3330 (RW)
0xa7: frame_vm_group_bin_19400 (RW)
0xa8: frame_vm_group_bin_12219 (RW)
0xa9: frame_vm_group_bin_5129 (RW)
0xa: frame_vm_group_bin_2931 (RW)
0xaa: frame_vm_group_bin_21225 (RW)
0xab: frame_vm_group_bin_14048 (RW)
0xac: frame_vm_group_bin_6857 (RW)
0xad: frame_vm_group_bin_23062 (RW)
0xae: frame_vm_group_bin_15879 (RW)
0xaf: frame_vm_group_bin_8688 (RW)
0xb0: frame_vm_group_bin_1499 (RW)
0xb1: frame_vm_group_bin_17639 (RW)
0xb2: frame_vm_group_bin_10510 (RW)
0xb3: frame_vm_group_bin_3363 (RW)
0xb4: frame_vm_group_bin_19432 (RW)
0xb5: frame_vm_group_bin_12251 (RW)
0xb6: frame_vm_group_bin_5162 (RW)
0xb7: frame_vm_group_bin_21258 (RW)
0xb8: frame_vm_group_bin_14081 (RW)
0xb9: frame_vm_group_bin_6882 (RW)
0xb: frame_vm_group_bin_19001 (RW)
0xba: frame_vm_group_bin_23096 (RW)
0xbb: frame_vm_group_bin_15913 (RW)
0xbc: frame_vm_group_bin_8722 (RW)
0xbd: frame_vm_group_bin_1533 (RW)
0xbe: frame_vm_group_bin_17673 (RW)
0xbf: frame_vm_group_bin_10543 (RW)
0xc0: frame_vm_group_bin_3394 (RW)
0xc1: frame_vm_group_bin_19463 (RW)
0xc2: frame_vm_group_bin_12285 (RW)
0xc3: frame_vm_group_bin_5196 (RW)
0xc4: frame_vm_group_bin_21292 (RW)
0xc5: frame_vm_group_bin_14115 (RW)
0xc6: frame_vm_group_bin_6906 (RW)
0xc7: frame_vm_group_bin_23129 (RW)
0xc8: frame_vm_group_bin_15946 (RW)
0xc9: frame_vm_group_bin_8755 (RW)
0xc: frame_vm_group_bin_11857 (RW)
0xca: frame_vm_group_bin_1566 (RW)
0xcb: frame_vm_group_bin_17701 (RW)
0xcc: frame_vm_group_bin_10576 (RW)
0xcd: frame_vm_group_bin_3418 (RW)
0xce: frame_vm_group_bin_19496 (RW)
0xcf: frame_vm_group_bin_12318 (RW)
0xd0: frame_vm_group_bin_5229 (RW)
0xd1: frame_vm_group_bin_21324 (RW)
0xd2: frame_vm_group_bin_14148 (RW)
0xd3: frame_vm_group_bin_6936 (RW)
0xd4: frame_vm_group_bin_23161 (RW)
0xd5: frame_vm_group_bin_15979 (RW)
0xd6: frame_vm_group_bin_8788 (RW)
0xd7: frame_vm_group_bin_1599 (RW)
0xd8: frame_vm_group_bin_17726 (RW)
0xd9: frame_vm_group_bin_10609 (RW)
0xd: frame_vm_group_bin_4732 (RW)
0xda: frame_vm_group_bin_3441 (RW)
0xdb: frame_vm_group_bin_19530 (RW)
0xdd: frame_vm_group_bin_5263 (RW)
0xe0: frame_vm_group_bin_6968 (RW)
0xe3: frame_vm_group_bin_8822 (RW)
0xe6: frame_vm_group_bin_10643 (RW)
0xe7: frame_vm_group_bin_3466 (RW)
0xe8: frame_vm_group_bin_19563 (RW)
0xe9: frame_vm_group_bin_12384 (RW)
0xe: frame_vm_group_bin_20851 (RW)
0xec: frame_vm_group_bin_14214 (RW)
0xed: frame_vm_group_bin_7001 (RW)
0xee: frame_vm_group_bin_23218 (RW)
0xef: frame_vm_group_bin_16048 (RW)
0xf2: frame_vm_group_bin_17784 (RW)
0xf3: frame_vm_group_bin_10674 (RW)
0xf4: frame_vm_group_bin_3492 (RW)
0xf5: frame_vm_group_bin_19597 (RW)
0xf: frame_vm_group_bin_13656 (RW)
}
pwm_obj_7_0_control_9_tcb {
cspace: pwm_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pwm_obj_group_bin_0305 (RW)
vspace: pwm_obj_group_bin_pd
}
pwm_obj_7_0_fault_handler_15_0000_tcb {
cspace: pwm_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pwm_obj_group_bin_0283 (RW)
vspace: pwm_obj_group_bin_pd
}
pwm_obj_7_i2c0_int_8_0000_tcb {
cspace: pwm_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pwm_obj_group_bin_0015 (RW)
vspace: pwm_obj_group_bin_pd
}
pwm_obj_7_pwm_3_0000_tcb {
cspace: pwm_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pwm_obj_group_bin_0061 (RW)
vspace: pwm_obj_group_bin_pd
}
pwm_obj_7_signal_6_0000_tcb {
cspace: pwm_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pwm_obj_group_bin_0286 (RW)
vspace: pwm_obj_group_bin_pd
}
pwm_obj_7_timer_update_12_0000_tcb {
cspace: pwm_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_pwm_obj_group_bin_0196 (RW)
vspace: pwm_obj_group_bin_pd
}
pwm_obj_cnode {
0x10: pwm_obj_pre_init_ep (RW)
0x11: pwm_obj_interface_init_ep (RW)
0x12: pwm_obj_post_init_ep (RW)
0x13: i2c0_irq_ntfn (R)
0x14: i2c0_irq_irq
0x15: pwm_sig_notification_0 (R)
0x16: pwm_sig_handoff_0 (RW)
0x17: pwm_sig_lock_0 (RW)
0x18: pwm_timer_notification_0 (R)
0x19: pwm_timer_handoff_0 (RW)
0x1: pwm_obj_set_motors (RW)
0x1a: pwm_timer_lock_0 (RW)
0x1b: fd_pwm.vm_pwm_ep (RW)
0x1c: pwm_obj_cnode (guard: 0, guard_size: 27)
0x2: pwm_obj_sig (RW)
0x3: pwm_obj_bus_sem (RW)
0x4: pwm_obj_7_0_control_9_tcb
0x5: pwm_obj_fault_ep (RWX, badge: 4)
0x6: pwm_obj_7_i2c0_int_8_0000_tcb
0x7: pwm_obj_fault_ep (RWX, badge: 6)
0x8: pwm_obj_7_signal_6_0000_tcb
0x9: pwm_obj_fault_ep (RWX, badge: 8)
0xa: pwm_obj_7_timer_update_12_0000_tcb
0xb: pwm_obj_fault_ep (RWX, badge: 10)
0xc: pwm_obj_7_pwm_3_0000_tcb
0xd: pwm_obj_fault_ep (RWX, badge: 12)
0xe: pwm_obj_7_0_fault_handler_15_0000_tcb
0xf: pwm_obj_fault_ep (RWX)
}
pwm_obj_group_bin_pd {
0x0: pt_pwm_obj_group_bin_0000
0x1: pt_pwm_obj_group_bin_0259
}
spi1_irq_irq {
0x0: spi1_irq_ntfn (R)
}
spi_obj_7_0_control_9_tcb {
cspace: spi_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_spi_obj_group_bin_0131 (RW)
vspace: spi_obj_group_bin_pd
}
spi_obj_7_0_fault_handler_15_0000_tcb {
cspace: spi_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_spi_obj_group_bin_0087 (RW)
vspace: spi_obj_group_bin_pd
}
spi_obj_7_spi1_int_8_0000_tcb {
cspace: spi_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_spi_obj_group_bin_0025 (RW)
vspace: spi_obj_group_bin_pd
}
spi_obj_7_spi_3_0000_tcb {
cspace: spi_obj_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_spi_obj_group_bin_0234 (RW)
vspace: spi_obj_group_bin_pd
}
spi_obj_cnode {
0x10: spi_clk_ep (WX, badge: 0)
0x11: can_spi_ep (RW)
0x12: spi_obj_cnode (guard: 0, guard_size: 27)
0x1: spi_obj_bus_sem (RW)
0x2: spi_obj_7_0_control_9_tcb
0x3: spi_obj_fault_ep (RWX, badge: 2)
0x4: spi_obj_7_spi1_int_8_0000_tcb
0x5: spi_obj_fault_ep (RWX, badge: 4)
0x6: spi_obj_7_spi_3_0000_tcb
0x7: spi_obj_fault_ep (RWX, badge: 6)
0x8: spi_obj_7_0_fault_handler_15_0000_tcb
0x9: spi_obj_fault_ep (RWX)
0xa: spi_obj_pre_init_ep (RW)
0xb: spi_obj_interface_init_ep (RW)
0xc: spi_obj_post_init_ep (RW)
0xd: spi1_irq_ntfn (R)
0xe: spi1_irq_irq
0xf: spi_gpio_ep (WX, badge: 0)
}
spi_obj_group_bin_pd {
0x0: pt_spi_obj_group_bin_0000
0x1: pt_spi_obj_group_bin_0247
}
timer_irq_irq {
0x0: timer_irq_ntfn (R)
}
timer_obj_9_0_control_9_tcb {
cspace: timer_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_timer_obj_group_bin_0084 (RW)
vspace: timer_obj_group_bin_pd
}
timer_obj_9_0_fault_handler_15_0000_tcb {
cspace: timer_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_timer_obj_group_bin_0179 (RW)
vspace: timer_obj_group_bin_pd
}
timer_obj_9_irq_3_0000_tcb {
cspace: timer_obj_cnode (guard: 0, guard_size: 28)
ipc_buffer_slot: frame_timer_obj_group_bin_0083 (RW)
vspace: timer_obj_group_bin_pd
}
timer_obj_cnode {
0x1: timer_obj_9_0_control_9_tcb
0x2: timer_obj_fault_ep (RWX, badge: 1)
0x3: timer_obj_9_irq_3_0000_tcb
0x4: timer_obj_fault_ep (RWX, badge: 3)
0x5: timer_obj_9_0_fault_handler_15_0000_tcb
0x6: timer_obj_fault_ep (RWX)
0x7: timer_obj_pre_init_ep (RW)
0x8: timer_obj_interface_init_ep (RW)
0x9: timer_obj_post_init_ep (RW)
0xa: pwm_timer_notification_0 (W)
0xb: timer_irq_ntfn (R)
0xc: timer_irq_irq
}
timer_obj_group_bin_pd {
0x0: pt_timer_obj_group_bin_0000
0x1: pt_timer_obj_group_bin_0235
}
uart_gcs_8_0_control_9_tcb {
cspace: uart_gcs_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_uart_gcs_group_bin_0026 (RW)
vspace: uart_gcs_group_bin_pd
}
uart_gcs_8_0_fault_handler_15_0000_tcb {
cspace: uart_gcs_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_uart_gcs_group_bin_0087 (RW)
vspace: uart_gcs_group_bin_pd
}
uart_gcs_8_interrupt_9_0000_tcb {
cspace: uart_gcs_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_uart_gcs_group_bin_0233 (RW)
vspace: uart_gcs_group_bin_pd
}
uart_gcs_8_uart_4_0000_tcb {
cspace: uart_gcs_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_uart_gcs_group_bin_0088 (RW)
vspace: uart_gcs_group_bin_pd
}
uart_gcs_cnode {
0x10: uart_inf_ep (RW)
0x11: uart_gcs_cnode (guard: 0, guard_size: 27)
0x13: gcs_recv_inf.px4_recv_inf_ep (WX, badge: 0)
0x1: uart_gcs_read_sem (RW)
0x2: uart_gcs_write_sem (RW)
0x3: uart_gcs_8_0_control_9_tcb
0x4: uart_gcs_fault_ep (RWX, badge: 3)
0x5: uart_gcs_8_interrupt_9_0000_tcb
0x6: uart_gcs_fault_ep (RWX, badge: 5)
0x7: uart_gcs_8_uart_4_0000_tcb
0x8: uart_gcs_fault_ep (RWX, badge: 7)
0x9: uart_gcs_8_0_fault_handler_15_0000_tcb
0xa: uart_gcs_fault_ep (RWX)
0xb: uart_gcs_pre_init_ep (RW)
0xc: uart_gcs_interface_init_ep (RW)
0xd: uart_gcs_post_init_ep (RW)
0xe: uartbase_irq_ntfn (R)
0xf: uartbase_irq_irq
}
uart_gcs_group_bin_pd {
0x0: pt_uart_gcs_group_bin_0000
0x1: pt_uart_gcs_group_bin_0246
}
uart_px4_8_0_control_9_tcb {
cspace: uart_px4_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_uart_px4_group_bin_0026 (RW)
vspace: uart_px4_group_bin_pd
}
uart_px4_8_0_fault_handler_15_0000_tcb {
cspace: uart_px4_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_uart_px4_group_bin_0087 (RW)
vspace: uart_px4_group_bin_pd
}
uart_px4_8_interrupt_9_0000_tcb {
cspace: uart_px4_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_uart_px4_group_bin_0233 (RW)
vspace: uart_px4_group_bin_pd
}
uart_px4_8_uart_4_0000_tcb {
cspace: uart_px4_cnode (guard: 0, guard_size: 27)
ipc_buffer_slot: frame_uart_px4_group_bin_0088 (RW)
vspace: uart_px4_group_bin_pd
}
uart_px4_cnode {
0x10: uartpx4_inf_ep (RW)
0x11: uart_px4_cnode (guard: 0, guard_size: 27)
0x13: gcs_recv_inf.px4_recv_inf_ep (WX, badge: 1)
0x1: uart_px4_read_sem (RW)
0x2: uart_px4_write_sem (RW)
0x3: uart_px4_8_0_control_9_tcb
0x4: uart_px4_fault_ep (RWX, badge: 3)
0x5: uart_px4_8_interrupt_9_0000_tcb
0x6: uart_px4_fault_ep (RWX, badge: 5)
0x7: uart_px4_8_uart_4_0000_tcb
0x8: uart_px4_fault_ep (RWX, badge: 7)
0x9: uart_px4_8_0_fault_handler_15_0000_tcb
0xa: uart_px4_fault_ep (RWX)
0xb: uart_px4_pre_init_ep (RW)
0xc: uart_px4_interface_init_ep (RW)
0xd: uart_px4_post_init_ep (RW)
0xe: uartpx4_irq_ntfn (R)
0xf: uartpx4_irq_irq
}
uart_px4_group_bin_pd {
0x0: pt_uart_px4_group_bin_0000
0x1: pt_uart_px4_group_bin_0246
}
uartbase_irq_irq {
0x0: uartbase_irq_ntfn (R)
}
uartpx4_irq_irq {
0x0: uartpx4_irq_ntfn (R)
}
vm_2_0_control_9_tcb {
cspace: vm_cnode (guard: 0, guard_size: 9)
ipc_buffer_slot: frame_vm_group_bin_8822 (RW)
vspace: vm_group_bin_pd
}
vm_2_0_fault_handler_15_0000_tcb {
cspace: vm_cnode (guard: 0, guard_size: 9)
ipc_buffer_slot: frame_vm_group_bin_5263 (RW)
vspace: vm_group_bin_pd
}
vm_2_restart_event_13_0000_tcb {
cspace: vm_cnode (guard: 0, guard_size: 9)
ipc_buffer_slot: frame_vm_group_bin_6968 (RW)
vspace: vm_group_bin_pd
}
vm_asid_pool {

}
vm_cnode {
0x10: vm_group_bin_pd
0x11: vm_simple_untyped_24_pool_0
0x12: vm_simple_untyped_24_pool_1
0x13: vm_simple_untyped_24_pool_2
0x14: vm_simple_untyped_24_pool_3
0x15: vm_simple_untyped_24_pool_4
0x16: vm_simple_untyped_24_pool_5
0x17: vm_simple_untyped_24_pool_6
0x18: vm_simple_untyped_24_pool_7
0x19: vm_simple_untyped_24_pool_8
0x1: vm_vm_sem (RW)
0x1a: vm_simple_untyped_24_pool_9
0x1b: vm_mmio_frame_268500992 (RW)
0x1c: vm_mmio_frame_268566528 (RW)
0x1d: vm_mmio_frame_322961408 (RW)
0x1e: vm_mmio_frame_268517376 (RW)
0x1f: vm_untyped_cap_268435456
0x20: vm_untyped_cap_273178624
0x21: vm_untyped_cap_314703872
0x22: vm_untyped_cap_268697600
0x23: vm_untyped_cap_268701696
0x24: vm_untyped_cap_268705792
0x25: vm_untyped_cap_268709888
0x26: vm_untyped_cap_268713984
0x27: vm_untyped_cap_268763136
0x28: vm_untyped_cap_268632064
0x29: vm_untyped_cap_268664832
0x2: vm_2_0_control_9_tcb
0x2a: vm_untyped_cap_268550144
0x2b: vm_untyped_cap_268533760
0x2c: vm_untyped_cap_303104000
0x2d: vm_untyped_cap_303235072
0x2e: vm_untyped_cap_304087040
0x2f: vm_untyped_cap_304218112
0x30: vm_untyped_cap_1073741824
0x31: vm_asid_pool
0x32: vm_irq_notification_obj (R)
0x33: vm_irq_27
0x34: vm_irq_85
0x35: vm_irq_107
0x36: vm_irq_109
0x37: vm_irq_103
0x3: vm_fault_ep (RWX, badge: 2)
0x4: vm_2_restart_event_13_0000_tcb
0x5: vm_fault_ep (RWX, badge: 4)
0x6: vm_2_0_fault_handler_15_0000_tcb
0x7: vm_fault_ep (RWX)
0x8: vm_pre_init_ep (RW)
0x9: vm_interface_init_ep (RW)
0xa: vm_post_init_ep (RW)
0xb: restart_vm_notification_0 (R)
0xc: restart_vm_handoff_0 (RW)
0xd: restart_vm_lock_0 (RW)
0xe: fd_pwm.vm_pwm_ep (WX, badge: 1)
0xf: vm_cnode (guard: 0, guard_size: 9)
}
vm_group_bin_pd {
0x0: pt_vm_group_bin_0000
0x10: pt_vm_group_bin_0006
0x11: pt_vm_group_bin_0044
0x12: pt_vm_group_bin_0065
0x13: pt_vm_group_bin_0031
0x14: pt_vm_group_bin_0117
0x15: pt_vm_group_bin_0051
0x16: pt_vm_group_bin_0014
0x17: pt_vm_group_bin_0167
0x18: pt_vm_group_bin_0004
0x19: pt_vm_group_bin_0033
0x1: pt_vm_group_bin_0063
0x1a: pt_vm_group_bin_0134
0x1b: pt_vm_group_bin_0022
0x1c: pt_vm_group_bin_0016
0x1d: pt_vm_group_bin_0008
0x1e: pt_vm_group_bin_0176
0x1f: pt_vm_group_bin_0035
0x20: pt_vm_group_bin_0054
0x21: pt_vm_group_bin_0328
0x22: pt_vm_group_bin_0018
0x23: pt_vm_group_bin_0010
0x24: pt_vm_group_bin_0037
0x25: pt_vm_group_bin_0060
0x26: pt_vm_group_bin_0024
0x27: pt_vm_group_bin_0020
0x28: pt_vm_group_bin_0210
0x29: pt_vm_group_bin_0012
0x2: pt_vm_group_bin_0028
0x2a: pt_vm_group_bin_0039
0x2b: pt_vm_group_bin_0403
0x2c: pt_vm_group_bin_0026
0x2d: pt_vm_group_bin_1120
0x3: pt_vm_group_bin_0220
0x4: pt_vm_group_bin_0002
0x5: pt_vm_group_bin_0099
0x6: pt_vm_group_bin_0380
0x7: pt_vm_group_bin_0196
0x8: pt_vm_group_bin_0071
0x9: pt_vm_group_bin_0272
0xa: pt_vm_group_bin_0079
0xb: pt_vm_group_bin_0239
0xc: pt_vm_group_bin_0123
0xd: pt_vm_group_bin_0203
0xe: pt_vm_group_bin_0115
0xf: pt_vm_group_bin_0107
}
vm_irq_103 {
0x0: vm_irq_notification_obj (R)
}
vm_irq_107 {
0x0: vm_irq_notification_obj (R)
}
vm_irq_109 {
0x0: vm_irq_notification_obj (R)
}
vm_irq_27 {
0x0: vm_irq_notification_obj (R)
}
vm_irq_85 {
0x0: vm_irq_notification_obj (R)
}
}

irq maps {
101: spi1_irq_irq
103: vm_irq_103
107: vm_irq_107
109: vm_irq_109
27: vm_irq_27
58: gpio_grp26_irq_irq
60: gpio_grp28_irq_irq
63: gpio_grp31_irq_irq
64: gpio_xint16_31_irq_irq
72: timer_irq_irq
84: uartpx4_irq_irq
85: vm_irq_85
86: uartbase_irq_irq
88: i2c0_irq_irq
}